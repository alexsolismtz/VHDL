library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY ROM_LUT_test64kx32 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END ROM_LUT_test64kx32;


architecture bijeibural of ROM_LUT_test64kx32 is
type RomType is array (natural range <>) of std_logic_vector(31 downto 0);
signal ROM : RomType(0 to 65535) := (

x"86936CA3",
x"86B46CC8",
x"86AB6CCB",
x"86776CA7",
x"861B6C61",
x"85A06BFA",
x"85096B7C",
x"84636AED",
x"83B86A59",
x"831369C9",
x"827C6949",
x"81FA68E1",
x"81946894",
x"814C6865",
x"81216852",
x"810D6856",
x"810A686C",
x"810E6889",
x"811468AB",
x"811368CC",
x"810468ED",
x"80E66910",
x"80B86934",
x"807D695C",
x"80356989",
x"7FE369B4",
x"7F8A69D9",
x"7F2A69EC",
x"7EC269E2",
x"7E5369B0",
x"7DDB694E",
x"7D5868BB",
x"7CCF67FD",
x"7C416720",
x"7BB46634",
x"7B2B654E",
x"7AAD647D",
x"7A3563D5",
x"79C46358",
x"79516307",
x"78CC62D8",
x"782762B7",
x"77526290",
x"763C624E",
x"74DF61E0",
x"733A613F",
x"7155606C",
x"6F485F70",
x"6D335E63",
x"6B3A5D5D",
x"69875C7E",
x"683E5BE0",
x"677D5B95",
x"67545BA9",
x"67C55C1C",
x"68C25CE3",
x"6A325DE9",
x"6BF05F14",
x"6DD16049",
x"6FAD616D",
x"715F626A",
x"72D16334",
x"73F463C4",
x"74C86418",
x"7559643B",
x"75BA6439",
x"76036421",
x"764B6401",
x"76AD63E8",
x"773763DD",
x"77F663EC",
x"78F06417",
x"7A24645D",
x"7B8764BE",
x"7D116535",
x"7EB265BE",
x"8058664E",
x"81EF66E0",
x"8366676D",
x"84AA67EF",
x"85AB685E",
x"865D68B7",
x"86BB68FC",
x"86C6692E",
x"868A6954",
x"86166976",
x"858669A3",
x"84F969E3",
x"84906A42",
x"846A6ACB",
x"84A16B7C",
x"85456C58",
x"865C6D55",
x"87DC6E69",
x"89B16F82",
x"8BC0708F",
x"8DE6717E",
x"8FFE7241",
x"91EA72D0",
x"93917325",
x"94E47344",
x"95DF7339",
x"96867312",
x"96E972E1",
x"971A72B9",
x"972B72A9",
x"973272BE",
x"973872FF",
x"9748736A",
x"976073F5",
x"977D7496",
x"97977537",
x"97A775C7",
x"97A47631",
x"978D766A",
x"97607665",
x"97227625",
x"96DD75AC",
x"9695750B",
x"96577451",
x"96277396",
x"960872EC",
x"95FC7266",
x"95FC7212",
x"960871F5",
x"961A7212",
x"962E725F",
x"964872D4",
x"96697361",
x"969A73F8",
x"96E3748B",
x"974F750D",
x"97E3757B",
x"98A275D1",
x"998B760F",
x"9A92763A",
x"9BAB7655",
x"9CBF7667",
x"9DB87671",
x"9E807677",
x"9F037677",
x"9F33766E",
x"9F0A765B",
x"9E857639",
x"9DAC7602",
x"9C8B75B7",
x"9B327557",
x"99B674E2",
x"982B745E",
x"96A273D0",
x"952F7340",
x"93E172B6",
x"92C9723B",
x"91EF71D8",
x"915A7195",
x"91117170",
x"9115716E",
x"915F718A",
x"91E771BE",
x"929F7200",
x"93747245",
x"944D7282",
x"951872A9",
x"95B972B3",
x"96217299",
x"963D7258",
x"960871EF",
x"9579715F",
x"949170AB",
x"934F6FD5",
x"91B26ED9",
x"8FB56DB5",
x"8D536C65",
x"8A816ADE",
x"8734691B",
x"8362671A",
x"7F0764D8",
x"7A2E625F",
x"74EA5FBC",
x"6F635D0A",
x"69CA5A63",
x"645E57E9",
x"5F5F55BA",
x"5B1153F4",
x"57AB52AC",
x"555151EB",
x"541651B0",
x"53F151F0",
x"54C45293",
x"565F537F",
x"58835495",
x"5AF155B6",
x"5D6656CA",
x"5FB157C0",
x"61AB588E",
x"63425930",
x"647659AC",
x"65575A0D",
x"65FF5A5C",
x"668F5AA5",
x"67255AF4",
x"67DF5B4D",
x"68CE5BB3",
x"69F95C26",
x"6B5B5CA1",
x"6CE95D21",
x"6E8C5D9E",
x"702D5E15",
x"71B45E84",
x"730E5EE9",
x"742B5F42",
x"75065F92",
x"759E5FDC",
x"75FC6021",
x"762B6063",
x"763B60A5",
x"763B60E9",
x"76376131",
x"763A617C",
x"764861CB",
x"7663621F",
x"76896279",
x"76B562D5",
x"76E66334",
x"771A6391",
x"775263ED",
x"77936446",
x"77E36498",
x"784C64E2",
x"78D16523",
x"7977655B",
x"7A3E6589",
x"7B2365B1",
x"7C1B65D5",
x"7D1D65F7",
x"7E16661B",
x"7EFC6645",
x"7FBF6675",
x"805866AD",
x"80C166ED",
x"80F66734",
x"80FA6780",
x"80D167CC",
x"80806813",
x"800D6851",
x"7F7C687D",
x"7ED36893",
x"7E14688D",
x"7D456869",
x"7C686827",
x"7B8067C9",
x"7A966752",
x"79AB66C9",
x"78CB6638",
x"77F665A4",
x"77326514",
x"76816490",
x"75E66418",
x"755F63AE",
x"74E86350",
x"747F62FC",
x"742062AB",
x"73C8625D",
x"7373620E",
x"732061C1",
x"72CC6174",
x"7279612D",
x"722460EE",
x"71CF60BB",
x"717A6094",
x"71276077",
x"70D5605F",
x"708A6043",
x"7046601D",
x"70115FE4",
x"6FED5F94",
x"6FDF5F2C",
x"6FE85EB1",
x"70095E2C",
x"70415DAC",
x"708D5D42",
x"70E85CFB",
x"714B5CE9",
x"71AE5D0E",
x"720C5D71",
x"725D5E0A",
x"72A05ECC",
x"72D55FA9",
x"72FD608D",
x"731D6168",
x"733B622B",
x"735C62CF",
x"7387634F",
x"73C263AE",
x"740D63F2",
x"746A6423",
x"74D66446",
x"754F6465",
x"75C9647F",
x"763E6491",
x"76A06497",
x"76DC6486",
x"76E36455",
x"76A063FA",
x"75FF6370",
x"74EC62AF",
x"735B61B8",
x"71426090",
x"6EA75F39",
x"6B945DC1",
x"68235C2F",
x"647A5A94",
x"60CA58FB",
x"5D455775",
x"5A29560C",
x"57A754D1",
x"55EE53D1",
x"551D5315",
x"554252A8",
x"565B528E",
x"584E52CE",
x"5AF85366",
x"5E245450",
x"619D5585",
x"652856FA",
x"6891589B",
x"6BAD5A59",
x"6E5C5C1F",
x"708A5DD7",
x"72355F70",
x"736360D5",
x"742161F9",
x"748662D0",
x"74A76358",
x"749A6391",
x"74736381",
x"743F6338",
x"740A62C4",
x"73D56239",
x"73A461AD",
x"73766132",
x"734760D9",
x"731660AB",
x"72E260AB",
x"72AB60D8",
x"72776128",
x"724C6191",
x"72346207",
x"7238627D",
x"726662ED",
x"72C86356",
x"736663BC",
x"7445642A",
x"756664A7",
x"76BF6544",
x"78466603",
x"79E866EB",
x"7B8D67F2",
x"7D23690C",
x"7E916A27",
x"7FCE6B2B",
x"80CE6C06",
x"81946CA6",
x"822D6D03",
x"82A76D1E",
x"831A6D06",
x"839E6CCB",
x"84446C87",
x"85186C51",
x"86206C3E",
x"87526C5B",
x"889F6CA8",
x"89F06D23",
x"8B2C6DBA",
x"8C3C6E5B",
x"8D106EF3",
x"8D9C6F70",
x"8DE36FCA",
x"8DEF6FF9",
x"8DD07002",
x"8D9C6FEF",
x"8D676FCA",
x"8D416F9D",
x"8D326F73",
x"8D396F51",
x"8D526F35",
x"8D696F1C",
x"8D6F6EFE",
x"8D4F6ED5",
x"8CFB6E9A",
x"8C6A6E4D",
x"8B986DEE",
x"8A8D6D80",
x"89536D0F",
x"87FD6CA0",
x"869E6C3B",
x"85496BE6",
x"84106BA3",
x"82FE6B70",
x"821E6B4B",
x"81726B2E",
x"80F66B10",
x"80A56AED",
x"80766ABE",
x"805D6A82",
x"80516A34",
x"804169D8",
x"8028696D",
x"7FFD68FC",
x"7FBA6883",
x"7F5B6809",
x"7EE36791",
x"7E536721",
x"7DB166BB",
x"7D00665E",
x"7C48660A",
x"7B8D65C1",
x"7AD5657D",
x"7A20653C",
x"797064FC",
x"78C564B5",
x"781E646A",
x"777A6417",
x"76D963BE",
x"763A6362",
x"75A06307",
x"750D62B1",
x"74836263",
x"74006221",
x"738361E9",
x"730661B7",
x"727F6181",
x"71E16141",
x"711E60EC",
x"702A6077",
x"6EFA5FDC",
x"6D895F1A",
x"6BD95E31",
x"69F75D2C",
x"67F85C18",
x"65F55B05",
x"640F5A0A",
x"626B5936",
x"6126589C",
x"605C5843",
x"60205833",
x"60795867",
x"616458D7",
x"62D15978",
x"64AA5A3C",
x"66D25B14",
x"69285BF3",
x"6B905CD2",
x"6DEC5DAB",
x"70285E83",
x"72385F5C",
x"7419603E",
x"75CF6131",
x"77656239",
x"78ED635D",
x"7A79649A",
x"7C1665E9",
x"7DCF6741",
x"7FAC6899",
x"81A869E1",
x"83BC6B10",
x"85D96C1D",
x"87F26D04",
x"89F66DC4",
x"8BDC6E62",
x"8DA26EE8",
x"8F4D6F61",
x"90E76FD8",
x"9283705C",
x"943270F9",
x"960D71B9",
x"981D72A0",
x"9A6D73B3",
x"9CFA74F1",
x"9FB87657",
x"A29277E0",
x"A5707982",
x"A8337B34",
x"AAC67CEB",
x"AD0E7E99",
x"AEFF802F",
x"B09881A2",
x"B1DC82E1",
x"B2DA83E6",
x"B3A884A7",
x"B45C8523",
x"B50F8560",
x"B5D98566",
x"B6C78542",
x"B7E08505",
x"B92384C2",
x"BA858487",
x"BBF4845E",
x"BD56844D",
x"BE918453",
x"BF8C8468",
x"C0378485",
x"C08884A3",
x"C08584B9",
x"C03D84C9",
x"BFCC84D7",
x"BF5784F4",
x"BF05852C",
x"BEFC8597",
x"BF5B8642",
x"C0378736",
x"C1918876",
x"C35D89F4",
x"C5848B9D",
x"C7E08D50",
x"CA4C8EF1",
x"CCA29060",
x"CEC69186",
x"D0A29253",
x"D23292C8",
x"D37692EF",
x"D48092D9",
x"D56092A0",
x"D623925D",
x"D6DA9224",
x"D7889200",
x"D82691F4",
x"D8AC91FA",
x"D9039203",
x"D9189200",
x"D8D491DF",
x"D8279196",
x"D705911B",
x"D56B9074",
x"D35E8FA8",
x"D0ED8EC3",
x"CE278DD8",
x"CB2C8CF4",
x"C8138C27",
x"C5048B7B",
x"C21B8AFA",
x"BF7B8AA7",
x"BD498A84",
x"BB9E8A94",
x"BA918AD9",
x"BA2D8B4F",
x"BA778BF6",
x"BB5E8CC5",
x"BCC78DB2",
x"BE888EAA",
x"C06D8F96",
x"C23A905C",
x"C3BA90E2",
x"C4B79110",
x"C50E90D5",
x"C4A8902B",
x"C3828F16",
x"C1AC8DA4",
x"BF418BEC",
x"BC688A0B",
x"B943881B",
x"B5F18635",
x"B2878466",
x"AF0782AD",
x"AB6A8107",
x"A7987F5D",
x"A37A7D9F",
x"9EF87BB3",
x"9A0A7989",
x"94B2771C",
x"8F0E7471",
x"894E7199",
x"83B26EB3",
x"7E896BE2",
x"7A1E694E",
x"76B5671A",
x"74806562",
x"73966438",
x"73F263A4",
x"7575639F",
x"77EB641D",
x"7B116509",
x"7EA7664C",
x"826967D6",
x"86256991",
x"89C16B75",
x"8D2E6D79",
x"90776F9A",
x"93B571DA",
x"97067437",
x"9A8B76B7",
x"9E637956",
x"A29B7C11",
x"A7397EE0",
x"AC3281B9",
x"B1708491",
x"B6D38757",
x"BC3A8A00",
x"C17C8C7A",
x"C67B8EB8",
x"CB1890B1",
x"CF40925C",
x"D2E893BA",
x"D61094CC",
x"D8BC959D",
x"DAF99637",
x"DCD596AD",
x"DE64970D",
x"DFB3976C",
x"E0D397D4",
x"E1C8984C",
x"E29A98D8",
x"E347996E",
x"E3C89A03",
x"E4169A89",
x"E4269AEF",
x"E3F59B26",
x"E37F9B26",
x"E2CB9AEE",
x"E1E49A85",
x"E0DA99F9",
x"DFC4995E",
x"DEBC98CA",
x"DDD89851",
x"DD2F9809",
x"DCCE97F9",
x"DCC0982A",
x"DD039897",
x"DD8F9937",
x"DE5099F9",
x"DF2C9ACB",
x"E0089B99",
x"E0C39C4E",
x"E13D9CD8",
x"E15E9D2A",
x"E1109D3D",
x"E04B9D0A",
x"DF109C99",
x"DD719BF1",
x"DB899B20",
x"D97F9A3E",
x"D7839961",
x"D5C3989F",
x"D46C9810",
x"D3A397C4",
x"D37997C5",
x"D3F49813",
x"D4FC98A3",
x"D66E9961",
x"D8139A2E",
x"D9AF9AEC",
x"DAFF9B78",
x"DBC89BB3",
x"DBE29B8A",
x"DB339AF2",
x"D9BD99EE",
x"D7989893",
x"D4F296FD",
x"D20C9555",
x"CF2D93C2",
x"CC9A926F",
x"CA909179",
x"C93A90F6",
x"C8AD90E9",
x"C8E29147",
x"C9C091F7",
x"CB1592D8",
x"CCA793C2",
x"CE3D948E",
x"CF9D9520",
x"D0A39563",
x"D13C9559",
x"D16A950C",
x"D1449493",
x"D0EF9410",
x"D09993A5",
x"D06A9370",
x"D0829382",
x"D0EE93DE",
x"D1A99479",
x"D29C953A",
x"D39D95FC",
x"D482969B",
x"D51D96F6",
x"D54D96F5",
x"D4FF968C",
x"D43695C7",
x"D30694B8",
x"D18E9382",
x"CFF19245",
x"CE4A9122",
x"CCA9902E",
x"CB048F69",
x"C93A8EC6",
x"C7198E27",
x"C4638D62",
x"C0D38C46",
x"BC388AAC",
x"B6778873",
x"AF948591",
x"A7BD820C",
x"9F407E08",
x"968A79B2",
x"8E147547",
x"865D7108",
x"7FD36D31",
x"7AC769F5",
x"77686773",
x"75BB65BC",
x"75A164CC",
x"76DB6490",
x"791464E9",
x"7BF065B1",
x"7F1866C5",
x"82416801",
x"8535694C",
x"87D86A93",
x"8A1F6BCA",
x"8C176CEE",
x"8DD36E00",
x"8F6D6F08",
x"90FD700A",
x"9291710D",
x"94327215",
x"95DA7320",
x"9780742F",
x"9911753A",
x"9A7A763E",
x"9BAC7731",
x"9C9C780D",
x"9D4B78CB",
x"9DBB7965",
x"9DFD79DA",
x"9E257A29",
x"9E4A7A56",
x"9E817A68",
x"9EDE7A65",
x"9F6A7A58",
x"A0297A49",
x"A1147A3E",
x"A21C7A40",
x"A32C7A51",
x"A42E7A6F",
x"A5047A9B",
x"A5997ACA",
x"A5E17AF9",
x"A5D07B1E",
x"A56C7B2F",
x"A4BB7B29",
x"A3D57B05",
x"A2CF7AC6",
x"A1C67A6E",
x"A0D77A06",
x"A01B799C",
x"9FA4793C",
x"9F7B78F5",
x"9FA878D7",
x"A02278E7",
x"A0DC7929",
x"A1C0799B",
x"A2B97A2F",
x"A3AB7AD4",
x"A47B7B78",
x"A5177C02",
x"A56C7C61",
x"A56E7C82",
x"A51F7C5E",
x"A4827BF4",
x"A3A57B4B",
x"A29A7A72",
x"A175797E",
x"A0547883",
x"9F52779C",
x"9E8776DE",
x"9E0B765B",
x"9DF47625",
x"9E4D7643",
x"9F1D76B7",
x"A0637783",
x"A21578A0",
x"A4257A05",
x"A67B7BA3",
x"A9007D6B",
x"AB997F50",
x"AE338143",
x"B0C08336",
x"B3328521",
x"B58986FB",
x"B7CA88C0",
x"B9FB8A70",
x"BC268C06",
x"BE518D81",
x"C07F8EDD",
x"C2A99016",
x"C4C49120",
x"C6BD91F2",
x"C87F9284",
x"C9F892CF",
x"CB1592D3",
x"CBCD9297",
x"CC1F9225",
x"CC139190",
x"CBB790EC",
x"CB22904F",
x"CA688FCB",
x"C99B8F6A",
x"C8C78F2E",
x"C7F58F10",
x"C71F8F00",
x"C63A8EE6",
x"C5368EA8",
x"C4018E32",
x"C28B8D6F",
x"C0C78C56",
x"BEB78AEA",
x"BC608938",
x"B9D48756",
x"B72D8560",
x"B4898378",
x"B20581BF",
x"AFB8804C",
x"ADAE7F2F",
x"ABE37E6B",
x"AA3F7DEF",
x"A89B7DA0",
x"A6C07D59",
x"A4767CE5",
x"A17D7C15",
x"9DA97ABA",
x"98E078B3",
x"932175F2",
x"8C90727F",
x"856D6E79",
x"7E116A16",
x"76E6659E",
x"705C615F",
x"6AD45DA7",
x"66A05AB8",
x"63EC58C3",
x"62C557DC",
x"631657FE",
x"64A45907",
x"67245AC0",
x"6A3F5CEA",
x"6D9D5F3C",
x"70EF6174",
x"73FA6362",
x"769764E0",
x"78B565E3",
x"7A536672",
x"7B8466A0",
x"7C5C6687",
x"7CF6664C",
x"7D6C6609",
x"7DCE65D6",
x"7E2B65C1",
x"7E8965CC",
x"7EEC65F9",
x"7F4F663B",
x"7FAF6689",
x"800966D5",
x"80556717",
x"80916749",
x"80BB6768",
x"80D16776",
x"80D26776",
x"80C2676D",
x"80A76760",
x"80866758",
x"80676753",
x"80566759",
x"805D6768",
x"8081677F",
x"80CB679A",
x"813867B8",
x"81C867D6",
x"827467EF",
x"83326803",
x"83F76813",
x"84B86826",
x"856A683F",
x"8607686C",
x"868D68B4",
x"86FC6920",
x"875869B7",
x"87AB6A79",
x"87FC6B63",
x"88556C6B",
x"88BE6D82",
x"893E6E94",
x"89DA6F90",
x"8A937062",
x"8B6970FF",
x"8C59715C",
x"8D5D717B",
x"8E717161",
x"8F8D7117",
x"90A770B0",
x"91B4703D",
x"92AA6FCB",
x"937E6F6B",
x"94286F21",
x"949F6EF2",
x"94DD6EDB",
x"94DF6ED5",
x"94A56EDB",
x"94346EE1",
x"93946EDF",
x"92D26ED4",
x"91F96EBB",
x"91186E99",
x"903E6E6E",
x"8F766E43",
x"8EC86E1C",
x"8E3B6E00",
x"8DCF6DF3",
x"8D836DF6",
x"8D4F6E06",
x"8D2E6E20",
x"8D176E3A",
x"8D016E4F",
x"8CE66E58",
x"8CBF6E4F",
x"8C8A6E31",
x"8C466DFD",
x"8BF36DBB",
x"8B916D6E",
x"8B256D21",
x"8AAF6CDC",
x"8A356CA6",
x"89B76C84",
x"89376C7A",
x"88B86C86",
x"883E6C9E",
x"87C86CBF",
x"875C6CDF",
x"86F76CF6",
x"869D6CFD",
x"864B6CF0",
x"85FD6CD1",
x"85B46CA0",
x"85696C61",
x"85186C1C",
x"84C16BD4",
x"84626B92",
x"83FF6B58",
x"839A6B28",
x"833E6B07",
x"82F26AF5",
x"82BE6AF0",
x"82A76AF9",
x"82AF6B0D",
x"82D26B28",
x"83016B45",
x"832E6B59",
x"833B6B59",
x"830E6B3A",
x"828B6AEC",
x"81976A65",
x"801D6999",
x"7E146886",
x"7B806730",
x"786F659E",
x"74FD63E2",
x"71566211",
x"6DAB6046",
x"6A2E5E9B",
x"67175D28",
x"64925C00",
x"62C45B2F",
x"61C55ABC",
x"619D5AA4",
x"62455AE1",
x"63A65B67",
x"659D5C25",
x"68035D0D",
x"6AAA5E0E",
x"6D635F1E",
x"7009602F",
x"7277613C",
x"7496623C",
x"7656632A",
x"77B26401",
x"78AE64C1",
x"79536562",
x"79B265E5",
x"79DD6648",
x"79E9668E",
x"79E666BB",
x"79E866D2",
x"79FA66DB",
x"7A2766DC",
x"7A7366DE",
x"7ADB66E0",
x"7B5B66E9",
x"7BE666F9",
x"7C72670D",
x"7CEF6727",
x"7D526741",
x"7D94675C",
x"7DB16776",
x"7DAB6790",
x"7D8D67AB",
x"7D6067CB",
x"7D3867EF",
x"7D236819",
x"7D2B6845",
x"7D5E6872",
x"7DB8689A",
x"7E3A68B7",
x"7ED668C2",
x"7F8168BA",
x"802D689A",
x"80CB6866",
x"81526820",
x"81BC67D1",
x"820B677D",
x"8242672E",
x"826966EC",
x"828466BB",
x"829B66A0",
x"82B2669A",
x"82C866AD",
x"82D966D3",
x"82DF670E",
x"82D26756",
x"82AE67A8",
x"826A6801",
x"82096859",
x"818B68AB",
x"80F768F2",
x"80586928",
x"7FB7694B",
x"7F21695C",
x"7EA2695B",
x"7E446951",
x"7E0B6942",
x"7DFD693C",
x"7E1A6949",
x"7E5C696F",
x"7EBF69B4",
x"7F3A6A19",
x"7FC46A97",
x"80516B24",
x"80D66BB4",
x"814F6C33",
x"81B26C93",
x"81FC6CC5",
x"822B6CC1",
x"82436C82",
x"824B6C0D",
x"82456B6D",
x"823B6AB2",
x"823469F0",
x"8237693B",
x"824368A6",
x"825F683E",
x"82816809",
x"82AA6806",
x"82CE682D",
x"82E8686D",
x"82ED68B4",
x"82DC68EC",
x"82AE6903",
x"826568EC",
x"820668A3",
x"81976828",
x"8122678A",
x"80B266DB",
x"80516632",
x"800365A7",
x"7FD1654C",
x"7FB76532",
x"7FB26559",
x"7FBB65BE",
x"7FC86653",
x"7FD16704",
x"7FCB67BB",
x"7FB16862",
x"7F8068E9",
x"7F3B6944",
x"7EE0696D",
x"7E756965",
x"7DF76930",
x"7D6568D2",
x"7CB4684C",
x"7BD5679E",
x"7AB866C4",
x"794C65B4",
x"77806465",
x"754B62D0",
x"72AE60F6",
x"6FB75EDD",
x"6C825C98",
x"69315A43",
x"65F357FD",
x"62FB55ED",
x"60765438",
x"5E8D52F8",
x"5D595243",
x"5CE8521F",
x"5D335287",
x"5E295367",
x"5FA954A2",
x"618C5618",
x"63A657A5",
x"65CF592B",
x"67E55A92",
x"69CA5BC9",
x"6B6D5CC9",
x"6CC85D92",
x"6DDC5E2E",
x"6EB15EA5",
x"6F555F08",
x"6FD65F64",
x"70465FC6",
x"70B46037",
x"712D60BE",
x"71BA615D",
x"72656218",
x"732E62E9",
x"741463CB",
x"751364B8",
x"762065A4",
x"77306684",
x"7834674E",
x"791E67F2",
x"79E06869",
x"7A6F68AA",
x"7AC468B0",
x"7ADE687C",
x"7AC16811",
x"7A77677A",
x"7A1166C5",
x"79A26601",
x"793C6544",
x"78F5649E",
x"78D96420",
x"78F363D5",
x"794863C8",
x"79D563FA",
x"7A936466",
x"7B746503",
x"7C6F65C1",
x"7D70668B",
x"7E6F6753",
x"7F5D6804",
x"8039688E",
x"80FE68EC",
x"81AE6919",
x"824E691A",
x"82E068FD",
x"837068D6",
x"840368B7",
x"84A068B5",
x"854B68E3",
x"8607694C",
x"86D669F5",
x"87B46AD8",
x"889D6BEB",
x"89876D17",
x"8A696E48",
x"8B356F65",
x"8BDF7058",
x"8C5D7112",
x"8CAA7189",
x"8CBF71BD",
x"8CA271B4",
x"8C59717C",
x"8BF17126",
x"8B7A70C3",
x"8B017061",
x"8A9A700A",
x"8A4E6FC7",
x"8A276F94",
x"8A296F70",
x"8A566F54",
x"8AA86F3A",
x"8B1D6F1C",
x"8BAC6EFA",
x"8C506ED9",
x"8D046EBD",
x"8DC26EAB",
x"8E836EB0",
x"8F3F6ECE",
x"8FEE6F08",
x"90886F5B",
x"91016FBE",
x"91527027",
x"9171708A",
x"915F70DC",
x"911B7113",
x"90AE712A",
x"90227121",
x"8F8A70FF",
x"8EF370CD",
x"8E6C7094",
x"8E007065",
x"8DB47045",
x"8D87703B",
x"8D737048",
x"8D6C7069",
x"8D667094",
x"8D5670C0",
x"8D3470E2",
x"8CFA70EF",
x"8CAC70DF",
x"8C4E70B1",
x"8BE97061",
x"8B856FF5",
x"8B2A6F72",
x"8AD66EDE",
x"8A816E3F",
x"8A1F6D9A",
x"899D6CEF",
x"88DF6C3A",
x"87CF6B76",
x"865B6A9C",
x"847669A4",
x"82236887",
x"7F6F6748",
x"7C7465E9",
x"79596476",
x"764662FE",
x"736C6197",
x"70F06053",
x"6EF35F46",
x"6D895E80",
x"6CB55E06",
x"6C725DD9",
x"6CAE5DF3",
x"6D515E46",
x"6E3E5EC3",
x"6F625F5C",
x"70AA6003",
x"720C60AF",
x"73876163",
x"75206221",
x"76E062F6",
x"78D163ED",
x"7AF66513",
x"7D586670",
x"7FF3680C",
x"82C469E1",
x"85C46BEB",
x"88ED6E1C",
x"8C387062",
x"8FA172B0",
x"932774F2",
x"96C5771C",
x"9A7A7923",
x"9E3C7B01",
x"A2037CB3",
x"A5BD7E3D",
x"A9597F9E",
x"ACBF80E0",
x"AFD98207",
x"B29B8319",
x"B4F58419",
x"B6E5850B",
x"B86B85F1",
x"B99286C9",
x"BA63878E",
x"BAEB883F",
x"BB3888D3",
x"BB518943",
x"BB3D898B",
x"BB0489A7",
x"BAA88994",
x"BA32895A",
x"B9AF8904",
x"B92D889F",
x"B8C3883F",
x"B88A87FB",
x"B89687E7",
x"B8FC8812",
x"B9C68887",
x"BAED8945",
x"BC658A3E",
x"BE0F8B5F",
x"BFC38C8A",
x"C1548D9E",
x"C2938E77",
x"C3588EFC",
x"C3898F17",
x"C31B8EC8",
x"C2158E17",
x"C0968D20",
x"BECA8C04",
x"BCE88AF3",
x"BB2C8A15",
x"B9D18995",
x"B904898F",
x"B8E68A11",
x"B97F8B1A",
x"BAC68C95",
x"BC9E8E65",
x"BED69060",
x"C1359259",
x"C3829423",
x"C5859599",
x"C712969D",
x"C80C9720",
x"C8689720",
x"C82F96A7",
x"C77895CC",
x"C66594AD",
x"C525936D",
x"C3E19232",
x"C2C4911D",
x"C1EB9048",
x"C16B8FC9",
x"C1498FA7",
x"C17B8FDB",
x"C1EA9052",
x"C27890F2",
x"C2FD9193",
x"C354920D",
x"C358923B",
x"C2F491FC",
x"C216913C",
x"C0C68FFA",
x"BF168E42",
x"BD2C8C35",
x"BB388A00",
x"B97087DA",
x"B80E85FE",
x"B73D84A1",
x"B72083E8",
x"B7C083ED",
x"B90B84AF",
x"BADC861B",
x"BCF58808",
x"BF0F8A42",
x"C0DE8C88",
x"C21D8EA0",
x"C29C9052",
x"C23F9176",
x"C10B91F6",
x"BF1F91D1",
x"BCAD9114",
x"B9F78FDB",
x"B7388E46",
x"B4A38C79",
x"B2538A8D",
x"B0498894",
x"AE648692",
x"AC71847E",
x"AA298246",
x"A7497FD6",
x"A3977D1B",
x"9EF47A06",
x"9966769D",
x"931472F1",
x"8C4C6F24",
x"85746B63",
x"7F0167E3",
x"796864DA",
x"75076277",
x"722460D8",
x"70DC6010",
x"7123601B",
x"72C960E9",
x"75846255",
x"78FA6438",
x"7CCE6665",
x"80AE68B1",
x"845F6AFD",
x"87BF6D30",
x"8AC56F3E",
x"8D807124",
x"900E72E5",
x"92947489",
x"95317619",
x"97FA7796",
x"9AF77905",
x"9E1B7A60",
x"A1527BA3",
x"A4767CC9",
x"A7677DCA",
x"AA057EA2",
x"AC387F53",
x"ADF57FE3",
x"AF408057",
x"B02580BA",
x"B0B98116",
x"B1158171",
x"B15081D4",
x"B1808243",
x"B1B582BC",
x"B1F78342",
x"B24C83CF",
x"B2B3845E",
x"B32C84EE",
x"B3B5857A",
x"B44E85FB",
x"B4FA8670",
x"B5BA86D7",
x"B694872E",
x"B7848774",
x"B88E87AC",
x"B9AC87DC",
x"BAD78805",
x"BC048833",
x"BD28886A",
x"BE3688AF",
x"BF25890A",
x"BFF0897A",
x"C09589FE",
x"C1188A93",
x"C17F8B2F",
x"C1D68BCF",
x"C2258C69",
x"C2748CF7",
x"C2C98D7B",
x"C3258DF4",
x"C3818E66",
x"C3D98ED6",
x"C4258F48",
x"C45E8FC2",
x"C4829042",
x"C49690C9",
x"C4A39151",
x"C4B691D3",
x"C4DE924B",
x"C52C92AE",
x"C5AC92FA",
x"C663932E",
x"C74E934E",
x"C864935E",
x"C9919365",
x"CAC1936F",
x"CBE19383",
x"CCE093AB",
x"CDB993EA",
x"CE6A9445",
x"CEFB94BA",
x"CF799544",
x"CFF795DB",
x"D07C9676",
x"D112970A",
x"D1B4978A",
x"D25A97EB",
x"D2EF9821",
x"D361982A",
x"D39A9802",
x"D39097AB",
x"D33D972E",
x"D2A79699",
x"D1E395F8",
x"D108955F",
x"D03994DE",
x"CF959484",
x"CF37945C",
x"CF36946D",
x"CF9994B8",
x"D0629538",
x"D18695E5",
x"D2EF96B1",
x"D4849790",
x"D627986F",
x"D7BA993E",
x"D91F99EE",
x"DA399A6E",
x"DAF19AB1",
x"DB379AB0",
x"DB039A65",
x"DA5199D1",
x"D92A98F8",
x"D79A97E5",
x"D5B496A5",
x"D38C9548",
x"D13493D9",
x"CEB39262",
x"CC0690E5",
x"C91B8F59",
x"C5D38DB1",
x"C2028BD3",
x"BD7A89A5",
x"B80F870D",
x"B1A583F1",
x"AA36804A",
x"A1D77C1E",
x"98BF777F",
x"8F457299",
x"85D66DA3",
x"7CEF68E1",
x"750C6495",
x"6E9A6101",
x"69EF5E57",
x"673D5CB6",
x"66895C26",
x"67B75C9A",
x"6A825DEA",
x"6E905FE6",
x"73786252",
x"78CC64F0",
x"7E2E678C",
x"834C69F9",
x"87EA6C20",
x"8BE76DF3",
x"8F346F75",
x"91D570B1",
x"93D971B7",
x"95577299",
x"966A735F",
x"97297415",
x"97A974B9",
x"97FD7548",
x"983375BD",
x"98567610",
x"986D7641",
x"987D7651",
x"98877646",
x"988B7626",
x"98887601",
x"987D75DC",
x"986675C3",
x"984375B9",
x"981A75BE",
x"97F075D1",
x"97CF75EC",
x"97C0760C",
x"97D0762F",
x"98077652",
x"98667678",
x"98ED76A5",
x"999576DB",
x"9A537720",
x"9B1B7772",
x"9BDF77D1",
x"9C987839",
x"9D40789F",
x"9DDA78FC",
x"9E6C7948",
x"9F00797E",
x"9FA47999",
x"A060799C",
x"A13C798F",
x"A239797C",
x"A355796E",
x"A4817975",
x"A5B3799C",
x"A6DC79EE",
x"A7EB7A6E",
x"A8D97B1F",
x"A9987BF7",
x"AA267CED",
x"AA807DEF",
x"AAA57EEB",
x"AA997FCD",
x"AA5E8088",
x"A9FB810B",
x"A9788151",
x"A8E1815D",
x"A8478136",
x"A7C380F0",
x"A76B809F",
x"A75D805D",
x"A7B08045",
x"A8748067",
x"A9B280D3",
x"AB61818B",
x"AD6A8287",
x"AFAB83B3",
x"B1F284F8",
x"B40F8638",
x"B5D08754",
x"B70B8831",
x"B7A988BE",
x"B7A388F0",
x"B70A88C9",
x"B5F88856",
x"B49887A7",
x"B31886D3",
x"B1A285EE",
x"B054850E",
x"AF42843D",
x"AE698381",
x"ADBC82DA",
x"AD218240",
x"AC7E81AC",
x"ABB68115",
x"AABC8075",
x"A98E7FCF",
x"A83A7F25",
x"A6E07E87",
x"A5A37DFF",
x"A4B17D9F",
x"A42C7D77",
x"A4317D8C",
x"A4C77DE5",
x"A5EA7E7E",
x"A77A7F46",
x"A94C802F",
x"AB2D8126",
x"ACE78212",
x"AE4782E1",
x"AF2C8384",
x"AF7E83F1",
x"AF3C8423",
x"AE6E841C",
x"AD2F83E0",
x"AB988372",
x"A9C282DC",
x"A7C3821B",
x"A5A3812D",
x"A35F8011",
x"A0E77EBD",
x"9E297D26",
x"9B0D7B46",
x"97817918",
x"938776A0",
x"8F2973E6",
x"8A8D7100",
x"85E36E06",
x"81706B1A",
x"7D7C6863",
x"7A4F6607",
x"782A642A",
x"773462E9",
x"7784625A",
x"79146284",
x"7BC26365",
x"7F5964EC",
x"839566FC",
x"882A6972",
x"8CC96C24",
x"91316EE6",
x"9529718F",
x"988E73FB",
x"9B4C760D",
x"9D5F77B6",
x"9ED378EE",
x"9FBE79B7",
x"A0387A22",
x"A05F7A3C",
x"A04A7A1C",
x"A01179D7",
x"9FBC797E",
x"9F54791D",
x"9ED978BC",
x"9E467858",
x"9D9577F1",
x"9CC2777C",
x"9BCC76F4",
x"9AB57652",
x"998A7597",
x"985874C7",
x"973573EF",
x"9639731F",
x"95797268",
x"950471E1",
x"94E37197",
x"95177195",
x"959271DB",
x"963D7264",
x"96FD731D",
x"97AF73F2",
x"983574C8",
x"98777586",
x"98667616",
x"97FE7667",
x"97497671",
x"96577636",
x"954575C1",
x"942C7525",
x"93287472",
x"924C73C4",
x"91A5732F",
x"913B72C4",
x"91087293",
x"910A72A0",
x"913572EB",
x"91817371",
x"91E77425",
x"926474F6",
x"92F375D5",
x"939076AD",
x"9435776C",
x"94DC77FF",
x"95747857",
x"95EE786B",
x"96397836",
x"964577BA",
x"96047703",
x"9573761F",
x"94977521",
x"937E7423",
x"9245733A",
x"9106727B",
x"8FE071F4",
x"8EF371AF",
x"8E5671AA",
x"8E1571E1",
x"8E387248",
x"8EB572D0",
x"8F7E7368",
x"90817402",
x"91A77496",
x"92D9751C",
x"94037596",
x"95147606",
x"96017672",
x"96C176DB",
x"974C7746",
x"97A177AC",
x"97B97808",
x"9798784E",
x"973C7874",
x"96B1786E",
x"95FE7836",
x"953877CB",
x"94777737",
x"93D9768D",
x"937B75E4",
x"937D7557",
x"93F97506",
x"94FB7508",
x"968D756C",
x"989E7639",
x"9B157764",
x"9DCC78D8",
x"A08B7A78",
x"A31E7C18",
x"A54A7D94",
x"A6E07EC6",
x"A7C07F91",
x"A7DC7FEA",
x"A7397FCD",
x"A5F77F4A",
x"A4407E7A",
x"A2507D77",
x"A05F7C64",
x"9E9D7B58",
x"9D297A6A",
x"9C117998",
x"9B3F78DD",
x"9A88781F",
x"99AE7741",
x"98647622",
x"966474A0",
x"937672A7",
x"8F74702D",
x"8A646D3B",
x"846A69EC",
x"7DCB6665",
x"76EB62DC",
x"703A5F87",
x"6A2B5C9C",
x"65275A46",
x"617958A6",
x"5F4F57C9",
x"5EB457AE",
x"5F8A5842",
x"619A5969",
x"64965AFB",
x"68265CD3",
x"6BF55EC8",
x"6FB760B8",
x"7334628B",
x"7645642E",
x"78DD6597",
x"7B0266C4",
x"7CC867B8",
x"7E4F687A",
x"7FB86917",
x"8127699C",
x"82B46A19",
x"84746A9E",
x"866F6B3A",
x"889F6BF8",
x"8AF96CE2",
x"8D676DFC",
x"8FCF6F43",
x"921470AB",
x"941B7226",
x"95CF739D",
x"971E74FB",
x"98037629",
x"987D7713",
x"989477AD",
x"985677F2",
x"97D577E7",
x"97247795",
x"9655770D",
x"95777665",
x"949575B0",
x"93B67502",
x"92DF7467",
x"921073E8",
x"914E738B",
x"909A734A",
x"8FF97320",
x"8F707308",
x"8F0672F8",
x"8EC372E8",
x"8EAF72D4",
x"8EC972B9",
x"8F157296",
x"8F8D726F",
x"90297248",
x"90E27223",
x"91A87206",
x"927071F0",
x"932B71E6",
x"93CF71E6",
x"945071EE",
x"94A771F8",
x"94CF7203",
x"94C67208",
x"948B7203",
x"942471F0",
x"939771CF",
x"92EF71A0",
x"92387166",
x"917E7124",
x"90D270E1",
x"904170A4",
x"8FD27072",
x"8F8D7051",
x"8F727041",
x"8F7C7043",
x"8FA17051",
x"8FD37066",
x"90047079",
x"90247080",
x"90257076",
x"8FFD7054",
x"8FA97017",
x"8F2B6FC4",
x"8E866F5C",
x"8DC66EEB",
x"8CF76E78",
x"8C246E0C",
x"8B586DB0",
x"8A9A6D68",
x"89ED6D35",
x"89506D16",
x"88BF6D04",
x"88346CF8",
x"87A76CE6",
x"87146CC7",
x"86766C93",
x"85CC6C44",
x"851E6BDC",
x"846F6B5B",
x"83C86AC7",
x"83356A2A",
x"82BE698C",
x"826868F6",
x"82376873",
x"8225680A",
x"822E67BC",
x"8242678E",
x"82556779",
x"82556779",
x"82326786",
x"81DF6794",
x"8153679A",
x"808D678E",
x"7F8E6769",
x"7E5F6725",
x"7D0B66C1",
x"7BA4663C",
x"7A32659E",
x"78C264EC",
x"7756642D",
x"75EA6366",
x"7478629B",
x"72ED61D0",
x"713B6100",
x"6F526027",
x"6D2B5F3F",
x"6AC85E43",
x"68345D32",
x"658A5C0D",
x"62F35AD7",
x"609D59A1",
x"5EB75877",
x"5D6F576E",
x"5CE8569C",
x"5D345614",
x"5E5555E3",
x"60355611",
x"62B2569F",
x"65995788",
x"68B158BD",
x"6BC45A2E",
x"6EA45BC2",
x"712D5D66",
x"73515F04",
x"750C608E",
x"766D61F9",
x"778E633C",
x"788E6459",
x"798C6553",
x"7AA06631",
x"7BDC66F9",
x"7D4667B5",
x"7EDB686C",
x"808D6921",
x"824869D8",
x"83F76A8D",
x"85866B3D",
x"86E06BE3",
x"87FC6C7A",
x"88D36CFD",
x"896C6D66",
x"89CE6DB5",
x"8A066DEC",
x"8A286E10",
x"8A466E26",
x"8A6F6E37",
x"8AAC6E48",
x"8B046E5E",
x"8B716E79",
x"8BEA6E94",
x"8C5C6EAA",
x"8CAE6EB0",
x"8CC86E99",
x"8C956E5B",
x"8C076DF0",
x"8B186D58",
x"89D56C97",
x"884F6BB8",
x"86A86ACF",
x"850B69ED",
x"83A2692B",
x"8294689B",
x"8200684B",
x"81F6683F",
x"82766877",
x"837068E9",
x"84C56983",
x"864C6A32",
x"87D66ADF",
x"89386B79",
x"8A4F6BF0",
x"8AFE6C3E",
x"8B3F6C5F",
x"8B146C5B",
x"8A8B6C3D",
x"89BC6C12",
x"88C56BE8",
x"87BF6BCC",
x"86C86BCC",
x"85F36BE9",
x"854C6C28",
x"84E06C86",
x"84B16CFD",
x"84C16D88",
x"850E6E1C",
x"859A6EB4",
x"86606F4B",
x"87606FDC",
x"88917066",
x"89EC70E6",
x"8B62715C",
x"8CE371C8",
x"8E5C7226",
x"8FB37275",
x"90D372AF",
x"91A872D1",
x"922172D5",
x"923572B9",
x"91E6727B",
x"91397217",
x"90417195",
x"8F1270F8",
x"8DCC7047",
x"8C8A6F8D",
x"8B6A6ED8",
x"8A846E33",
x"89E96DA9",
x"89A46D45",
x"89B16D0F",
x"8A096D08",
x"8A976D2E",
x"8B426D7A",
x"8BEA6DE2",
x"8C716E54",
x"8CBB6EBE",
x"8CAF6F0D",
x"8C3C6F30",
x"8B5C6F1C",
x"8A0E6EC8",
x"88636E37",
x"866A6D72",
x"84426C8A",
x"82066B93",
x"7FD86AA6",
x"7DD569D8",
x"7C14693E",
x"7AAA68E1",
x"799D68C1",
x"78ED68D5",
x"788D690A",
x"786B6945",
x"78696969",
x"78676958",
x"784668F9",
x"77E9683E",
x"77386723",
x"762865AF",
x"74BD63F9",
x"7300621D",
x"710E603E",
x"6F075E7D",
x"6D145CFA",
x"6B5E5BCC",
x"6A065B00",
x"692B5A98",
x"68E15A8E",
x"692B5AD3",
x"6A055B53",
x"6B5E5BFD",
x"6D215CBD",
x"6F345D8E",
x"717C5E67",
x"73DF5F4B",
x"764E6041",
x"78B86152",
x"7B1A6289",
x"7D7063E9",
x"7FBC6575",
x"82036728",
x"844868F9",
x"86916AD9",
x"88DF6CB7",
x"8B2E6E80",
x"8D777023",
x"8FB2718F",
x"91D072BB",
x"93C6739D",
x"95877436",
x"97077485",
x"98457492",
x"99437468",
x"9A0E7419",
x"9AB673B4",
x"9B527350",
x"9BF672FF",
x"9CB572D2",
x"9D9872D4",
x"9E997309",
x"9FA2736B",
x"A08D73EA",
x"A1267468",
x"A13674C7",
x"A08374E2",
x"9EDD749A",
x"9C2C73D5",
x"986D7288",
x"93BC70B4",
x"8E536E70",
x"887E6BE2",
x"829E6938",
x"7D1066A8",
x"782E6466",
x"743D629E",
x"7163616C",
x"6FAE60DD",
x"6F0960E9",
x"6F48617A",
x"7030626C",
x"717A6394",
x"72E864C5",
x"744165D8",
x"755E66AD",
x"762B6731",
x"76A4675F",
x"76D4673A",
x"76D166D5",
x"76B26644",
x"769365A3",
x"7683650B",
x"768F6494",
x"76B7644B",
x"76F56439",
x"7738645F",
x"776964B1",
x"776F651E",
x"77306590",
x"769765EC",
x"759A661D",
x"74386610",
x"728365BB",
x"709B6520",
x"6EB1644E",
x"6D02635F",
x"6BD26279",
x"6B6561C3",
x"6BF5616A",
x"6DA76190",
x"708A624C",
x"748D63AB",
x"798265A0",
x"7F1D6814",
x"85016ADE",
x"8AC66DCD",
x"900870A9",
x"94737343",
x"97C6756C",
x"99E3770B",
x"9ACC780F",
x"9AA47879",
x"999F7857",
x"980877C3",
x"962B76DA",
x"944D75BC",
x"92AA7485",
x"91627351",
x"9088722F",
x"901A7129",
x"90017045",
x"90256F88",
x"90646EEB",
x"90A56E70",
x"90D86E17",
x"90F36DDE",
x"90FB6DC8",
x"90FB6DD5",
x"91016E08",
x"911A6E59",
x"914C6EC4",
x"91946F3B",
x"91E06FAE",
x"92177006",
x"920E702E",
x"919B700F",
x"90906F93",
x"8EC56EA9",
x"8C216D4B",
x"88986B79",
x"8435693E",
x"7F1366B0",
x"796563EC",
x"736A6115",
x"6D6E5E53",
x"67BA5BCB",
x"6297599E",
x"5E4357E3",
x"5AE856AB",
x"58A155F7",
x"577355C2",
x"574F55F8",
x"58175684",
x"59A3574C",
x"5BC15835",
x"5E435928",
x"60FB5A14",
x"63C25AEE",
x"667C5BB1",
x"69135C5C",
x"6B765CF4",
x"6DA15D7D",
x"6F915DFC",
x"71485E76",
x"72C75EEA",
x"74135F5A",
x"75315FC5",
x"76276028",
x"76FC6081",
x"77B260D3",
x"7852611B",
x"78DB615D",
x"794E619B",
x"79A761D9",
x"79E36215",
x"79F96250",
x"79E06287",
x"799362B5",
x"790E62D6",
x"785362E4",
x"776962DC",
x"765F62BC",
x"75426287",
x"742B6242",
x"732B61F7",
x"725561B1",
x"71B7617E",
x"7158616A",
x"713A6181",
x"715961C8",
x"71AB6241",
x"722462E8",
x"72B563B1",
x"7353648D",
x"73F0656A",
x"74846635",
x"750766DB",
x"7576674B",
x"75CE677F",
x"760B6770",
x"76346724",
x"764566A4",
x"764465FD",
x"76326542",
x"76136483",
x"75EC63D0",
x"75BF6338",
x"759462C1",
x"756D6270",
x"754E6246",
x"753A623E",
x"75376253",
x"7545627E",
x"756C62B9",
x"75AD62FE",
x"76096349",
x"76816394",
x"771663E0",
x"77BF6427",
x"78766469",
x"792D64A4",
x"79D564D2",
x"7A5D64F0",
x"7AB764FA",
x"7AD564ED",
x"7AAF64C6",
x"7A496487",
x"79A8642F",
x"78E263C5",
x"780E6350",
x"774962DC",
x"76B16274",
x"76626229",
x"76706206",
x"76E8621A",
x"77C9626A",
x"790C62FD",
x"7A9863D0",
x"7C5664DC",
x"7E276611",
x"7FEA675C",
x"818468A6",
x"82DF69D9",
x"83EA6AE1",
x"849E6BAA",
x"84FD6C2B",
x"850A6C63",
x"84D06C54",
x"845D6C07",
x"83BF6B8D",
x"83066AF7",
x"823E6A56",
x"817369B7",
x"80B26927",
x"800468AB",
x"7F706845",
x"7EFA67F2",
x"7EA467AD",
x"7E6A676D",
x"7E48672E",
x"7E2E66E9",
x"7E106697",
x"7DD96634",
x"7D7765BC",
x"7CD6652D",
x"7BE86484",
x"7AA163C2",
x"790062E4",
x"770A61ED",
x"74C960E2",
x"72565FC8",
x"6FCA5EAB",
x"6D425D95",
x"6AE35C9B",
x"68CC5BCB",
x"671B5B33",
x"65EC5AE6",
x"65515AEB",
x"65545B46",
x"65F85BF7",
x"67375CF1",
x"69025E28",
x"6B3F5F88",
x"6DD560FE",
x"709D6274",
x"737363DA",
x"76346521",
x"78C16641",
x"7AFE6737",
x"7CDF6807",
x"7E5868B8",
x"7F706952",
x"803169DF",
x"80AE6A66",
x"81016AED",
x"81416B79",
x"81836C04",
x"81D96C90",
x"824F6D16",
x"82E86D8F",
x"839E6DF6",
x"846A6E48",
x"85416E82",
x"86116EA3",
x"86CF6EAB",
x"87706EA1",
x"87EC6E86",
x"883E6E5E",
x"88676E2D",
x"886A6DF5",
x"884B6DBA",
x"880D6D79",
x"87B76D34",
x"874D6CE9",
x"86DB6C99",
x"86656C44",
x"85F66BE9",
x"859D6B8D",
x"85636B35",
x"85586AE8",
x"85866AAD",
x"85F46A8F",
x"86A46A93",
x"87906AC2",
x"88AA6B1E",
x"89E06BA7",
x"8B1B6C57",
x"8C426D1E",
x"8D416DF2",
x"8E066EBF",
x"8E8B6F76",
x"8ED27008",
x"8EE3706B",
x"8ECF709C",
x"8EAA709D",
x"8E847076",
x"8E6D7035",
x"8E6C6FE6",
x"8E806F93",
x"8E9E6F44",
x"8EB76EFC",
x"8EB76EB5",
x"8E876E6C",
x"8E1B6E14",
x"8D676DA4",
x"8C6D6D16",
x"8B396C69",
x"89DF6BA4",
x"887C6AD4",
x"872C6A0A",
x"8614695E",
x"854E68E3",
x"84ED68AD",
x"850168C8",
x"858A693A",
x"868169FF",
x"87D26B09",
x"89646C47",
x"8B1A6DA0",
x"8CD06EF9",
x"8E6A7039",
x"8FC87148",
x"90D37216",
x"91807296",
x"91C572C5",
x"91A872A9",
x"9138724B",
x"908671BB",
x"8FAF7110",
x"8ED0705C",
x"8E066FB5",
x"8D6D6F2D",
x"8D186ED1",
x"8D186EA7",
x"8D716EB4",
x"8E226EF5",
x"8F1F6F62",
x"905A6FF3",
x"91BC709A",
x"932C714D",
x"949271FF",
x"95D272A4",
x"96D77334",
x"978D73A5",
x"97E373EE",
x"97D3740C",
x"975873FB",
x"967373B9",
x"952C7344",
x"939072A3",
x"91AC71D8",
x"8F8D70E9",
x"8D3E6FDE",
x"8AC66EBA",
x"88276D7F",
x"855C6C2D",
x"825D6ABF",
x"7F226931",
x"7BA4677A",
x"77E5659A",
x"73EC6390",
x"6FD56163",
x"6BC45F24",
x"67E85CEA",
x"647A5AD5",
x"61B35904",
x"5FC25799",
x"5ECE56B2",
x"5EE45660",
x"600256A8",
x"62095784",
x"64CD58E0",
x"680F5A9C",
x"6B8E5C95",
x"6F0D5EA2",
x"725860A1",
x"75476276",
x"77CC640D",
x"79E56560",
x"7BA16675",
x"7D196752",
x"7E66680A",
x"7FA268AE",
x"80E3694F",
x"823169F6",
x"838E6AAD",
x"84F76B75",
x"86656C4D",
x"87CF6D2D",
x"89326E12",
x"8A906EF6",
x"8BED6FD2",
x"8D5670A6",
x"8ED6716B",
x"90767221",
x"923B72CA",
x"94287364",
x"963573F1",
x"98567475",
x"9A7774F5",
x"9C887578",
x"9E777603",
x"A03376A0",
x"A1B37752",
x"A2F4781F",
x"A3F77903",
x"A4BF79F8",
x"A5567AF1",
x"A5C27BDE",
x"A60F7CAF",
x"A6437D50",
x"A6677DB5",
x"A6817DD9",
x"A69B7DBC",
x"A6BD7D6A",
x"A6F57CF2",
x"A74C7C6D",
x"A7CD7BEF",
x"A8827B92",
x"A96E7B61",
x"AA8C7B65",
x"ABD37B9F",
x"AD2F7C04",
x"AE8A7C86",
x"AFC57D16",
x"B0C97DA3",
x"B17B7E1E",
x"B1D07E7F",
x"B1C37EC9",
x"B15B7EFA",
x"B0AE7F1C",
x"AFD37F3A",
x"AEEB7F5D",
x"AE157F8A",
x"AD667FC0",
x"ACEB7FFC",
x"ACA68037",
x"AC8B8064",
x"AC858077",
x"AC7A8064",
x"AC4F8020",
x"ABED7FA9",
x"AB457EFE",
x"AA547E20",
x"A9227D19",
x"A7BF7BF4",
x"A6407ABC",
x"A4C0797F",
x"A352784A",
x"A205772A",
x"A0E17629",
x"9FE47550",
x"9F0A74A5",
x"9E45742C",
x"9D8B73E6",
x"9CD673D2",
x"9C1E73EC",
x"9B67742C",
x"9AB57485",
x"9A0D74EA",
x"9977754E",
x"98F675A2",
x"988775DB",
x"982775F2",
x"97CA75E1",
x"976675AC",
x"96F07555",
x"966074E8",
x"95AF7471",
x"94E373F9",
x"9403738C",
x"9318732F",
x"923272E1",
x"915F72A4",
x"90A97274",
x"901A7247",
x"8FB2721A",
x"8F6E71E9",
x"8F4971B4",
x"8F37717B",
x"8F297143",
x"8F12710F",
x"8EE070E1",
x"8E8470B7",
x"8DEA708A",
x"8D047051",
x"8BC46FF8",
x"8A1D6F6E",
x"880A6EA1",
x"858B6D88",
x"82AD6C1A",
x"7F7D6A5C",
x"7C1B685F",
x"78AD663C",
x"75596411",
x"72516204",
x"6FC16037",
x"6DD15ECB",
x"6CA05DD5",
x"6C425D64",
x"6CC15D7B",
x"6E175E12",
x"70315F1A",
x"72F5607E",
x"7644622B",
x"79F9640B",
x"7DF36610",
x"8214682E",
x"863F6A62",
x"8A626CA7",
x"8E6C6F00",
x"9253716C",
x"960E73E8",
x"9995766C",
x"9CE378EA",
x"9FEE7B50",
x"A2AE7D88",
x"A5157F78",
x"A71B810E",
x"A8B58235",
x"A9DC82E0",
x"AA8E830B",
x"AACA82BD",
x"AA988200",
x"AA0180E7",
x"A9157F8B",
x"A7E67E0B",
x"A68D7C7F",
x"A5237B05",
x"A3C579B7",
x"A28E78AC",
x"A19E77F5",
x"A10E77A0",
x"A0FA77B6",
x"A1717839",
x"A2827925",
x"A42C7A6E",
x"A6677C06",
x"A91F7DD7",
x"AC307FC3",
x"AF7581B3",
x"B2C2838A",
x"B5E7852F",
x"B8BD8691",
x"BB2687A5",
x"BD0F886D",
x"BE7788F0",
x"BF68893F",
x"BFFE896D",
x"C0578994",
x"C09589C5",
x"C0D68A10",
x"C1338A7D",
x"C1B68B0E",
x"C25D8BBB",
x"C31E8C79",
x"C3E38D36",
x"C4958DE7",
x"C51E8E7C",
x"C56F8EEC",
x"C5848F34",
x"C55E8F58",
x"C5108F5D",
x"C4AF8F4F",
x"C4518F35",
x"C4118F1B",
x"C3FB8F06",
x"C4198EF7",
x"C4678EEC",
x"C4DA8EE2",
x"C55B8ECE",
x"C5D48EAA",
x"C62C8E6C",
x"C64A8E10",
x"C6228D93",
x"C5AC8CF6",
x"C4EB8C3F",
x"C3ED8B76",
x"C2C48AA8",
x"C18C89E2",
x"C0608931",
x"BF5A88A2",
x"BE92883F",
x"BE1B880E",
x"BDFB8814",
x"BE35884C",
x"BEBF88B4",
x"BF85893F",
x"C07189E3",
x"C1688A91",
x"C24C8B3E",
x"C3078BD9",
x"C3858C5C",
x"C3C08CBE",
x"C3B48CFD",
x"C36D8D1A",
x"C2F98D1A",
x"C26D8D04",
x"C1D78CE2",
x"C1498CB9",
x"C0C38C91",
x"C0468C6A",
x"BFC38C42",
x"BF268C11",
x"BE5B8BCC",
x"BD4E8B67",
x"BBF08AD6",
x"BA378A0E",
x"B82F890A",
x"B5E487C8",
x"B36A864A",
x"B0D9849C",
x"AE4382C7",
x"ABAF80D7",
x"A9167ED3",
x"A6637CBD",
x"A3717A93",
x"A0147851",
x"9C2175EB",
x"97717355",
x"91F37088",
x"8BAB6D82",
x"84BC6A4B",
x"7D6266F5",
x"75F0639D",
x"6ECB6067",
x"68555D7D",
x"62EB5B04",
x"5ED4591C",
x"5C3A57DD",
x"5B2A574C",
x"5B895760",
x"5D245804",
x"5FB45915",
x"62E15A6B",
x"66595BDF",
x"69CF5D48",
x"6D075E8D",
x"6FDB5F9D",
x"72356076",
x"7417611D",
x"758D61A1",
x"76B16218",
x"77A06297",
x"7876632B",
x"794963E0",
x"7A2F64BA",
x"7B3165AF",
x"7C5066B7",
x"7D8D67C1",
x"7EDB68BE",
x"802D699C",
x"81726A51",
x"82956AD2",
x"838A6B1E",
x"843E6B3A",
x"84A86B2A",
x"84C56AFA",
x"84976AB8",
x"842B6A73",
x"83956A3A",
x"82EF6A1C",
x"82536A23",
x"81DD6A59",
x"81A56AC4",
x"81B96B61",
x"82236C2B",
x"82DA6D16",
x"83D66E10",
x"84FF6F08",
x"86396FE6",
x"876D709A",
x"88807112",
x"895D7145",
x"89FC7133",
x"8A5970E1",
x"8A7A705C",
x"8A6D6FB9",
x"8A436F0A",
x"8A0D6E69",
x"89DD6DE8",
x"89BF6D90",
x"89BB6D6C",
x"89CF6D78",
x"89FA6DAD",
x"8A346DFF",
x"8A736E62",
x"8AB26EC7",
x"8AED6F23",
x"8B276F70",
x"8B626FAD",
x"8BAA6FD7",
x"8C096FF3",
x"8C877008",
x"8D2C7017",
x"8DFA7029",
x"8EED703E",
x"8FF97057",
x"910D7070",
x"9215708A",
x"92FD70A1",
x"93AE70B1",
x"941870B9",
x"942F70B5",
x"93ED70A6",
x"93567089",
x"9274705F",
x"91597029",
x"90176FE6",
x"8EC96F9C",
x"8D846F4A",
x"8C606EF5",
x"8B6D6EA1",
x"8AB56E52",
x"8A3C6E0C",
x"8A006DCF",
x"89F96D9E",
x"8A156D76",
x"8A496D52",
x"8A866D30",
x"8ABB6D08",
x"8AE46CD8",
x"8AFE6C9D",
x"8B0A6C57",
x"8B116C0A",
x"8B1B6BBE",
x"8B326B79",
x"8B5D6B47",
x"8BA46B2E",
x"8C036B34",
x"8C746B5B",
x"8CF06BA1",
x"8D696C00",
x"8DD26C6D",
x"8E1E6CDC",
x"8E436D41",
x"8E3F6D8F",
x"8E0D6DBE",
x"8DB46DCB",
x"8D356DB4",
x"8C9A6D79",
x"8BE66D20",
x"8B1D6CAA",
x"8A396C1C",
x"89346B75",
x"87FD6AB0",
x"868369C7",
x"84B168B2",
x"82726768",
x"7FBA65E3",
x"7C846421",
x"78D66227",
x"74C76003",
x"70765DC6",
x"6C165B8D",
x"67DB5973",
x"64025795",
x"60C25611",
x"5E4B54F8",
x"5CC05459",
x"5C305436",
x"5C9A5489",
x"5DEB5547",
x"6002565D",
x"62AE57B9",
x"65C15945",
x"69065AED",
x"6C515CA7",
x"6F775E62",
x"725D6017",
x"74F361C1",
x"772B635A",
x"790964DE",
x"7A916646",
x"7BD16791",
x"7CD968BB",
x"7DBC69BF",
x"7E8E6AA0",
x"7F626B5F",
x"80466BFF",
x"81496C87",
x"826F6CFD",
x"83B56D68",
x"85156DCA",
x"867E6E23",
x"87E26E76",
x"89276EBF",
x"8A3E6EFC",
x"8B176F27",
x"8BAE6F41",
x"8C036F48",
x"8C1E6F40",
x"8C106F2D",
x"8BEC6F13",
x"8BC66EFA",
x"8BB26EE6",
x"8BBC6ED9",
x"8BEF6ED4",
x"8C466ED4",
x"8CC36ED7",
x"8D5C6ED8",
x"8E076ED7",
x"8EBC6ECF",
x"8F766EC8",
x"90316EC4",
x"90F16ECE",
x"91BB6EEF",
x"92976F34",
x"938B6FA7",
x"94A4704E",
x"95E3712B",
x"974D723D",
x"98E0737B",
x"9A9174D7",
x"9C56763E",
x"9E1B779D",
x"9FCF78DE",
x"A15C79EE",
x"A2AF7AC0",
x"A3BB7B4A",
x"A4767B8E",
x"A4DE7B91",
x"A4FA7B61",
x"A4D47B12",
x"A4817AB9",
x"A4117A6A",
x"A3987A37",
x"A3267A29",
x"A2C37A44",
x"A2707A84",
x"A22B7AD8",
x"A1E67B30",
x"A1987B78",
x"A1347B9C",
x"A0B07B8F",
x"A00F7B4B",
x"9F537AD0",
x"9E8B7A2C",
x"9DC8796E",
x"9D1E78AD",
x"9CA57801",
x"9C6A777B",
x"9C78772C",
x"9CCC7716",
x"9D5D7736",
x"9E177782",
x"9EDD77E8",
x"9F927856",
x"A01878B3",
x"A05278F1",
x"A02B7902",
x"9F9978E2",
x"9EA1788F",
x"9D4C7810",
x"9BB3776E",
x"99F976B7",
x"983F75F9",
x"96B17544",
x"956A74A1",
x"94877420",
x"941273C3",
x"940A7390",
x"945F7388",
x"94F373A5",
x"95A273DF",
x"9646742D",
x"96BB7482",
x"96DF74D0",
x"96A47509",
x"96047527",
x"95077520",
x"93BF74F1",
x"92457499",
x"90B1741A",
x"8F177378",
x"8D8172B6",
x"8BEF71D4",
x"8A5570D4",
x"88A26FB5",
x"86C16E76",
x"849D6D19",
x"822E6BA0",
x"7F726A14",
x"7C7C6884",
x"79666701",
x"765C659E",
x"738C6472",
x"7124638A",
x"6F5162F7",
x"6E3362BE",
x"6DDC62DC",
x"6E4F6349",
x"6F8063F4",
x"715864CB",
x"73B265BC",
x"766A66B4",
x"795967A7",
x"7C59688A",
x"7F51695B",
x"82256A1C",
x"84CC6ACF",
x"873E6B7A",
x"89796C24",
x"8B846CD2",
x"8D666D86",
x"8F256E41",
x"90CB6F03",
x"92596FC8",
x"93D5708D",
x"953B714D",
x"968A7202",
x"97BE72A6",
x"98D27339",
x"99C373B6",
x"9A91741F",
x"9B407479",
x"9BD674CB",
x"9C5F751D",
x"9CE37578",
x"9D7075E8",
x"9E117671",
x"9ECD7719",
x"9FA777DE",
x"A09B78B9",
x"A1AB79A3",
x"A2CD7A8F",
x"A3FD7B72",
x"A5397C44",
x"A6837D02",
x"A7DF7DAC",
x"A9557E47",
x"AAED7EE0",
x"ACB27F7E",
x"AEA5802F",
x"B0C380F8",
x"B2FF81DA",
x"B54682D0",
x"B77B83CC",
x"B98184BF",
x"BB39859B",
x"BC8B864D",
x"BD6586D2",
x"BDC38721",
x"BDAA8743",
x"BD2C8743",
x"BC638732",
x"BB6D871F",
x"BA6B8721",
x"B97C8742",
x"B8BA878A",
x"B83987FB",
x"B8078892",
x"B82B8946",
x"B8A98A0E",
x"B9828ADD",
x"BAB28BAC",
x"BC358C74",
x"BDFE8D2F",
x"C0028DDC",
x"C2328E79",
x"C4778F04",
x"C6BA8F7C",
x"C8E08FDD",
x"CACB9025",
x"CC67904E",
x"CD9C9052",
x"CE5E9032",
x"CEA78FEF",
x"CE798F8C",
x"CDDE8F0E",
x"CCE78E83",
x"CBA88DF4",
x"CA378D6D",
x"C8AD8CF7",
x"C71C8C9D",
x"C5948C62",
x"C4228C45",
x"C2CA8C45",
x"C1928C59",
x"C0778C77",
x"BF748C95",
x"BE848CAA",
x"BDA08CA8",
x"BCCA8C8D",
x"BBFF8C55",
x"BB468C01",
x"BAA38B98",
x"BA258B24",
x"B9CE8AAE",
x"B9A88A3F",
x"B9AF89E2",
x"B9D98998",
x"BA118962",
x"BA3F8939",
x"BA438915",
x"BA0288EE",
x"B96688B9",
x"B861886E",
x"B6FE880E",
x"B550879B",
x"B37D871E",
x"B1AF86A1",
x"B0148631",
x"AECC85D0",
x"ADE4857E",
x"AD50852F",
x"ACEB84CD",
x"AC718438",
x"AB95834D",
x"AA0181ED",
x"A7717FFC",
x"A3B37D6E",
x"9EBC7A46",
x"98A87699",
x"91BC7292",
x"8A5C6E65",
x"83036A52",
x"7C2E6696",
x"764F6369",
x"71BF60F7",
x"6EB45F5C",
x"6D3A5E9D",
x"6D375EAF",
x"6E755F78",
x"70A860D3",
x"737F6293",
x"76AA648B",
x"79E96693",
x"7D106889",
x"80076A55",
x"82C86BE8",
x"855D6D3D",
x"87D66E52",
x"8A466F34",
x"8CBB6FEC",
x"8F387089",
x"91BC7119",
x"943C71A9",
x"96A77245",
x"98E972F9",
x"9AF073C7",
x"9CAC74AF",
x"9E1A75AF",
x"9F3376C0",
x"A00477D7",
x"A09A78E8",
x"A10479EB",
x"A15A7AD3",
x"A1B37B96",
x"A2247C32",
x"A2BC7CA5",
x"A3857CED",
x"A4857D12",
x"A5B97D18",
x"A7157D06",
x"A88A7CE7",
x"AA027CC1",
x"AB6A7C9E",
x"ACAC7C86",
x"ADB67C81",
x"AE847C98",
x"AF0F7CD1",
x"AF637D32",
x"AF8A7DBF",
x"AF997E78",
x"AFA97F5B",
x"AFCD8064",
x"B0168187",
x"B08E82B5",
x"B13583E0",
x"B20084F6",
x"B2E185E7",
x"B3C286A7",
x"B489872C",
x"B5298777",
x"B58F878A",
x"B5BD876E",
x"B5B88736",
x"B59486EE",
x"B56886AC",
x"B554867E",
x"B5758671",
x"B5E0868B",
x"B6A086D0",
x"B7B9873B",
x"B91C87C2",
x"BAB6885D",
x"BC678900",
x"BE11899E",
x"BF988A2F",
x"C0E78AAE",
x"C1F48B17",
x"C2C08B69",
x"C3548BAA",
x"C3C78BDC",
x"C42D8C04",
x"C49E8C27",
x"C5298C48",
x"C5DA8C69",
x"C6AF8C8D",
x"C79F8CB2",
x"C8998CD9",
x"C9878CFB",
x"CA4E8D17",
x"CAD78D25",
x"CB0F8D21",
x"CAE48D00",
x"CA508CBE",
x"C9538C52",
x"C7F18BB8",
x"C6368AF0",
x"C43689FD",
x"C20888E9",
x"BFC487C0",
x"BD8B8699",
x"BB758588",
x"B9A384A5",
x"B82C8405",
x"B71E83B9",
x"B68283C9",
x"B6548436",
x"B68484F3",
x"B6F585EC",
x"B7858704",
x"B80A8818",
x"B85B8907",
x"B85789B1",
x"B7E489FB",
x"B6F789DA",
x"B58F894A",
x"B3BD8853",
x"B199870B",
x"AF42858A",
x"ACD483EC",
x"AA678249",
x"A80580B3",
x"A5AF7F35",
x"A3597DCA",
x"A0EB7C63",
x"9E4A7AEA",
x"9B5A7948",
x"98057768",
x"94457539",
x"901F72BA",
x"8BAC6FF6",
x"87176D06",
x"82906A10",
x"7E536741",
x"7A9764C5",
x"778E62C5",
x"75596160",
x"740C60A7",
x"73A36094",
x"740C6118",
x"75246214",
x"76C16362",
x"78B464D8",
x"7AD2664F",
x"7CF967AE",
x"7F0E68E2",
x"810769E5",
x"82E06ABE",
x"84A76B7C",
x"86656C31",
x"882A6CEE",
x"8A036DBE",
x"8BF96EAB",
x"8E0B6FB1",
x"903570CA",
x"926D71E6",
x"94A572FB",
x"96D273F8",
x"98EA74D8",
x"9AE77596",
x"9CCC7636",
x"9E9776C0",
x"A04D773E",
x"A1F077BC",
x"A380783E",
x"A4F478CD",
x"A6457965",
x"A7637A05",
x"A8437AA2",
x"A8D97B33",
x"A9257BB0",
x"A9307C16",
x"A90B7C63",
x"A8D77C9B",
x"A8B97CC6",
x"A8D97CEF",
x"A95D7D25",
x"AA647D71",
x"AC017DDE",
x"AE327E71",
x"B0EB7F2B",
x"B40F800A",
x"B77B8105",
x"BB018218",
x"BE788336",
x"C1BA8456",
x"C4AD8570",
x"C73C867E",
x"C95D877D",
x"CB0F886A",
x"CC578948",
x"CD3C8A15",
x"CDC68AD5",
x"CDFC8B87",
x"CDEB8C2E",
x"CD998CC6",
x"CD108D50",
x"CC5E8DC8",
x"CB8C8E2A",
x"CAA88E70",
x"C9BD8E98",
x"C8D48E9E",
x"C7F28E81",
x"C7188E42",
x"C6418DE3",
x"C5678D65",
x"C4848CCE",
x"C38E8C24",
x"C2878B6C",
x"C16E8AAB",
x"C04D89E7",
x"BF308928",
x"BE2A8871",
x"BD4A87C8",
x"BCA28732",
x"BC3C86B6",
x"BC1C8656",
x"BC428618",
x"BCA085FA",
x"BD2885FB",
x"BDC08617",
x"BE4F8643",
x"BEB38673",
x"BED38697",
x"BE9886A1",
x"BDEF8684",
x"BCD48638",
x"BB4C85B8",
x"B966850A",
x"B7428438",
x"B5098353",
x"B2ED8271",
x"B11B81A6",
x"AFC08104",
x"AF018098",
x"AEEB8064",
x"AF7F8064",
x"B0A5808A",
x"B23280BC",
x"B3ED80E4",
x"B59580E7",
x"B6ED80B3",
x"B7C28039",
x"B7F07F75",
x"B76B7E74",
x"B63F7D40",
x"B48B7BF4",
x"B27E7AAA",
x"B050797B",
x"AE33787C",
x"AC5277B9",
x"AABC7733",
x"A97376E2",
x"A86076B4",
x"A75A7693",
x"A62F7664",
x"A4A8760C",
x"A29A7575",
x"9FE47492",
x"9C82735C",
x"988771DA",
x"941B7019",
x"8F7A6E2E",
x"8AEA6C38",
x"86B56A54",
x"831868A1",
x"8048673C",
x"7E5D663C",
x"7D6265AE",
x"7D446595",
x"7DE365F0",
x"7F1466AE",
x"80A767BB",
x"826D68FC",
x"84446A55",
x"86116BAE",
x"87C86CF3",
x"896C6E16",
x"8B076F13",
x"8CAA6FEF",
x"8E6570B9",
x"904B717E",
x"92647255",
x"94B87350",
x"973F747B",
x"99F375DC",
x"9CC37774",
x"9FA27934",
x"A2807B0F",
x"A54D7CEF",
x"A8007EBD",
x"AA918064",
x"ACF881D6",
x"AF358305",
x"B14683EE",
x"B3268491",
x"B4D184F4",
x"B6428523",
x"B76E852C",
x"B850851F",
x"B8E0850A",
x"B91884F7",
x"B8FB84F4",
x"B88C8504",
x"B7D78529",
x"B6EE8563",
x"B5E985A8",
x"B4E185EE",
x"B3F4862C",
x"B33D8652",
x"B2D48656",
x"B2CF8631",
x"B33385DE",
x"B4078563",
x"B53F84C9",
x"B6CC8421",
x"B894837E",
x"BA7882F7",
x"BC5A829F",
x"BE18828A",
x"BF9882BC",
x"C0C3833C",
x"C18B8400",
x"C1EE84F7",
x"C1F1860E",
x"C19F872B",
x"C10B8832",
x"C049890A",
x"BF6D899E",
x"BE8889E2",
x"BDA689CD",
x"BCD08966",
x"BC0488B2",
x"BB4387C5",
x"BA8786B5",
x"B9CD8598",
x"B915848A",
x"B85E83A3",
x"B7B382FB",
x"B719829E",
x"B69F8297",
x"B65382E6",
x"B6408387",
x"B671846A",
x"B6EA857B",
x"B7AB86A4",
x"B8AC87C6",
x"B9E188CC",
x"BB36899D",
x"BC918A24",
x"BDD18A58",
x"BEDB8A32",
x"BF8E89B6",
x"BFCD88EC",
x"BF8287E3",
x"BEA586AE",
x"BD36855E",
x"BB42840E",
x"B8E782CD",
x"B64A81AF",
x"B39B80BD",
x"B10A8000",
x"AEC37F7B",
x"ACEA7F29",
x"AB947F02",
x"AAC57EFB",
x"AA717EFF",
x"AA7D7F04",
x"AAC27EF5",
x"AB157EC4",
x"AB4D7E6A",
x"AB477DDD",
x"AAEB7D22",
x"AA337C40",
x"A9267B44",
x"A7D47A3E",
x"A65C7943",
x"A4DA7864",
x"A36A77AF",
x"A21C7727",
x"A0F576CE",
x"9FED7696",
x"9EE77668",
x"9DC27627",
x"9C4D75B3",
x"9A5C74EA",
x"97C373B1",
x"946971F8",
x"90416FB9",
x"8B536D00",
x"85C169E6",
x"7FBE6691",
x"79916331",
x"73895FF3",
x"6DF55D08",
x"69205A9A",
x"654758C0",
x"628F578B",
x"610656FA",
x"60A45701",
x"61445787",
x"62B05871",
x"64A6599E",
x"66E25AEE",
x"69235C49",
x"6B355D98",
x"6CF35ECD",
x"6E4C5FE2",
x"6F4460CF",
x"6FEB6197",
x"7062623F",
x"70CC62C9",
x"7151633E",
x"720C63A3",
x"731163FC",
x"74696450",
x"760D64A7",
x"77EC6506",
x"79E9656F",
x"7BE965E5",
x"7DCC6668",
x"7F7966F7",
x"80DD678C",
x"81EF6820",
x"82AD68AA",
x"831E6920",
x"8352697A",
x"835969B2",
x"834869C7",
x"833169B8",
x"831F698C",
x"8321694C",
x"83376904",
x"836568C4",
x"83A56894",
x"83F3687F",
x"8446688A",
x"849A68B7",
x"84E668FF",
x"852B695C",
x"856569C5",
x"85986A31",
x"85CE6A97",
x"860D6AF5",
x"86626B48",
x"86D66B96",
x"87736BE1",
x"883F6C2E",
x"893B6C87",
x"8A5F6CEC",
x"8B9E6D5C",
x"8CE66DD2",
x"8E1E6E48",
x"8F316EB3",
x"90076F0C",
x"90936F4B",
x"90CC6F6F",
x"90B56F7A",
x"905A6F75",
x"8FD06F65",
x"8F316F59",
x"8E976F58",
x"8E1E6F6B",
x"8DD76F93",
x"8DD06FCE",
x"8E077016",
x"8E777064",
x"8F1070AD",
x"8FC170E9",
x"90747114",
x"911B712D",
x"91A97133",
x"9217712E",
x"92627123",
x"928B7117",
x"9298710F",
x"928D710A",
x"926D7106",
x"923970FE",
x"91F170E8",
x"919370BE",
x"911B707E",
x"90877020",
x"8FD86FAA",
x"8F0E6F20",
x"8E2F6E8A",
x"8D3C6DEF",
x"8C3F6D5C",
x"8B396CD5",
x"8A2F6C63",
x"89276C07",
x"88216BC4",
x"87256B99",
x"863B6B83",
x"856C6B86",
x"84C86BA0",
x"84606BD5",
x"84456C27",
x"84836C99",
x"85226D2A",
x"86226DD7",
x"87796E99",
x"890D6F62",
x"8AC27026",
x"8C7370D4",
x"8DFA715A",
x"8F3871AD",
x"901471C7",
x"907D71A4",
x"9074714E",
x"8FFE70CB",
x"8F2C702E",
x"8E116F83",
x"8CBC6ED8",
x"8B396E34",
x"898D6D96",
x"87B26CF8",
x"85A06C4E",
x"83486B8A",
x"80A56AA0",
x"7DB46983",
x"7A7E6832",
x"771D66B4",
x"73B2651B",
x"7069637D",
x"6D6F61F9",
x"6AF360A8",
x"69145FA5",
x"67E95F00",
x"67755EBD",
x"67AA5ED9",
x"686F5F42",
x"699C5FE2",
x"6B09609D",
x"6C91615A",
x"6E146204",
x"6F80628E",
x"70CB62F4",
x"71F96338",
x"73166366",
x"7434638B",
x"756363B9",
x"76B063FF",
x"78216466",
x"79B764F3",
x"7B6A65A7",
x"7D31667C",
x"7EFA6768",
x"80BB6860",
x"82696958",
x"83FD6A44",
x"857A6B1A",
x"86DF6BD1",
x"88356C62",
x"89836CCB",
x"8ACC6D0A",
x"8C116D21",
x"8D526D13",
x"8E866CE5",
x"8FA46CA1",
x"909F6C51",
x"916F6BFD",
x"92076BB1",
x"92666B76",
x"928A6B52",
x"927D6B4C",
x"924C6B68",
x"920D6BA4",
x"91D36C03",
x"91B66C86",
x"91CF6D2D",
x"922C6DF8",
x"92D96EE9",
x"93DD7002",
x"95327141",
x"96D072A1",
x"98A7741F",
x"9AA175A9",
x"9CA97734",
x"9EAB78AA",
x"A09279F9",
x"A2507B0F",
x"A3DD7BDB",
x"A5317C57",
x"A64D7C82",
x"A7327C63",
x"A7E67C0C",
x"A86D7B92",
x"A8C77B0F",
x"A8FB7A9D",
x"A9077A54",
x"A8E97A43",
x"A8A47A71",
x"A8367AE0",
x"A7A57B82",
x"A6FA7C49",
x"A63F7D20",
x"A5827DEF",
x"A4D67EA6",
x"A4497F33",
x"A3E97F91",
x"A3BB7FBD",
x"A3C37FBC",
x"A3FA7F98",
x"A4527F5B",
x"A4B67F0F",
x"A5147EBD",
x"A5537E64",
x"A5637E07",
x"A5367D9E",
x"A4C97D26",
x"A41C7C9B",
x"A33B7BF7",
x"A22F7B3A",
x"A10B7A68",
x"9FDD7986",
x"9EB278A0",
x"9D9277BC",
x"9C7E76E0",
x"9B777612",
x"9A777554",
x"997A74A5",
x"987B7400",
x"977B7365",
x"967C72D0",
x"9583723E",
x"949571B3",
x"93BC7130",
x"92FA70B7",
x"9250704F",
x"91BB6FF8",
x"91326FB3",
x"90AB6F7C",
x"901B6F4E",
x"8F7A6F27",
x"8EC86F02",
x"8E076EDB",
x"8D456EB4",
x"8C906E90",
x"8BFB6E72",
x"8B9A6E61",
x"8B706E5B",
x"8B806E5F",
x"8BB66E66",
x"8BF66E61",
x"8C156E3D",
x"8BE36DE3",
x"8B316D42",
x"89D56C47",
x"87B46AE9",
x"84C9692B",
x"812A6719",
x"7CFD64C9",
x"7881625C",
x"73FF5FF4",
x"6FC55DB9",
x"6C1A5BC9",
x"69385A3D",
x"67445925",
x"66475880",
x"66345847",
x"66EE586B",
x"683E58D6",
x"69F25973",
x"6BD25A2B",
x"6DAE5AEE",
x"6F635BB5",
x"70E15C7A",
x"721E5D41",
x"73255E0B",
x"74075EE3",
x"74D55FCD",
x"75A860CE",
x"769061E6",
x"779D6313",
x"78D26450",
x"7A356597",
x"7BBF66DF",
x"7D696821",
x"7F2A6954",
x"80F36A72",
x"82B96B76",
x"84736C5C",
x"86106D21",
x"878A6DC4",
x"88D96E45",
x"89F96EA7",
x"8AE76EEE",
x"8BA86F1D",
x"8C406F40",
x"8CB86F59",
x"8D156F70",
x"8D5F6F89",
x"8D9A6FA6",
x"8DC86FC4",
x"8DE66FDF",
x"8DF16FF2",
x"8DE66FF3",
x"8DBF6FDC",
x"8D7B6FAB",
x"8D206F5C",
x"8CB16EF5",
x"8C366E7A",
x"8BBE6DF6",
x"8B506D73",
x"8AF66CFC",
x"8AB16C96",
x"8A836C48",
x"8A626C14",
x"8A456BF6",
x"8A216BE8",
x"89E96BE6",
x"89976BE8",
x"89256BE9",
x"88976BE6",
x"87F76BDF",
x"87526BD9",
x"86B76BD5",
x"86386BDB",
x"85E26BEF",
x"85C16C16",
x"85D86C4F",
x"86286C9C",
x"86AF6CF6",
x"87606D5B",
x"88326DBE",
x"89176E1A",
x"8A006E65",
x"8AE06E96",
x"8BA76EAA",
x"8C466E9A",
x"8CB46E6B",
x"8CE26E1D",
x"8CCB6DBA",
x"8C6A6D4B",
x"8BC66CDB",
x"8AE76C78",
x"89E06C2E",
x"88C86C07",
x"87BC6C0A",
x"86D96C3A",
x"86366C93",
x"85E96D10",
x"85F66DA4",
x"865C6E3F",
x"87086ED1",
x"87E06F47",
x"88C26F8F",
x"89876F9C",
x"8A106F65",
x"8A416EE8",
x"8A0B6E26",
x"896F6D28",
x"88796C00",
x"873F6AC1",
x"85E56980",
x"848A6855",
x"834F6755",
x"824C6691",
x"81946616",
x"812765E6",
x"81006603",
x"810E6662",
x"813E66F5",
x"817767A8",
x"81A86869",
x"81BF6921",
x"81B569BC",
x"81866A2B",
x"81376A61",
x"80CC6A55",
x"80516A04",
x"7FC66975",
x"7F3268A7",
x"7E8E67A8",
x"7DD36683",
x"7CF36542",
x"7BE263F3",
x"7A91629F",
x"78FC6152",
x"771D600E",
x"75025EDC",
x"72B85DBF",
x"705F5CBC",
x"6E165BD5",
x"6C025B10",
x"6A485A73",
x"69095A04",
x"685C59CD",
x"685459D7",
x"68F05A28",
x"6A2D5AC5",
x"6BFA5BB1",
x"6E455CE9",
x"70F75E69",
x"73FA6028",
x"773B621B",
x"7AAB6435",
x"7E3C666C",
x"81E968B5",
x"85A76B04",
x"896D6D54",
x"8D316F9C",
x"90E371D5",
x"947373F9",
x"97CD7601",
x"9AE177E4",
x"9DA2799B",
x"A0037B1E",
x"A2017C68",
x"A3A47D75",
x"A4F07E47",
x"A5F67EDE",
x"A6C07F3F",
x"A75D7F70",
x"A7D27F74",
x"A81F7F50",
x"A8427F05",
x"A8307E95",
x"A7DD7DFC",
x"A73F7D3A",
x"A6507C53",
x"A5127B4A",
x"A38C7A2A",
x"A1D37902",
x"A00077E2",
x"9E2C76E0",
x"9C7A760C",
x"9B007575",
x"99CF7527",
x"98EE7523",
x"985D7564",
x"980D75DC",
x"97EA767E",
x"97E27733",
x"97E077E7",
x"97D87888",
x"97C57909",
x"97AB7962",
x"97957993",
x"9795799D",
x"97B87988",
x"9808795B",
x"988A7920",
x"993478E0",
x"99F178A0",
x"9AAB7862",
x"9B427829",
x"9B9C77F1",
x"9BA277B7",
x"9B4D777B",
x"9A9F7737",
x"99A976EA",
x"98887693",
x"975C7634",
x"964675D0",
x"95667567",
x"94CD7501",
x"948874A0",
x"9497744A",
x"94EF7403",
x"958373D2",
x"964373BB",
x"972473C6",
x"981773F4",
x"991B744B",
x"9A2B74CE",
x"9B48757C",
x"9C6E7652",
x"9D9A774B",
x"9EB9785B",
x"9FBE7974",
x"A08E7A85",
x"A1147B78",
x"A1397C39",
x"A0F07CB7",
x"A0357CE1",
x"9F0E7CAD",
x"9D917C1B",
x"9BD77B2C",
x"9A0579F1",
x"983F787B",
x"96A776E4",
x"9555754A",
x"945773C8",
x"93B47276",
x"93607168",
x"934870A7",
x"93527035",
x"93597009",
x"933E7012",
x"92E07039",
x"92287062",
x"91067076",
x"8F76705E",
x"8D7B700A",
x"8B2B6F76",
x"889F6EA3",
x"85F66D9C",
x"83526C70",
x"80D26B35",
x"7E9169FA",
x"7C9D68CE",
x"7AF967B8",
x"799866B8",
x"786665C4",
x"773F64CF",
x"75FF63C6",
x"747D629B",
x"72986142",
x"703B5FB3",
x"6D5C5DF7",
x"6A075C1A",
x"66565A32",
x"6272585D",
x"5E9256B8",
x"5AEB555D",
x"57BA5463",
x"552C53D4",
x"536853B3",
x"528053F5",
x"52785489",
x"53415556",
x"54BE5642",
x"56CA5735",
x"59375818",
x"5BD958E0",
x"5E8A5985",
x"61295A0B",
x"639D5A7A",
x"65D75ADD",
x"67D15B42",
x"698C5BB2",
x"6B0D5C35",
x"6C5B5CCF",
x"6D7C5D7A",
x"6E765E31",
x"6F4F5EEA",
x"700C5F9D",
x"70AE603C",
x"713C60C5",
x"71B86132",
x"72276187",
x"728A61C6",
x"72E661F4",
x"733D621B",
x"738C6241",
x"73D36266",
x"74106291",
x"744262BF",
x"746862ED",
x"7482631A",
x"74966341",
x"74A8635D",
x"74C26373",
x"74EC6380",
x"752B6387",
x"7584638E",
x"75F7639A",
x"767F63AD",
x"771363C9",
x"77AA63F2",
x"78346423",
x"78AA6458",
x"79006490",
x"793764C6",
x"794E64F9",
x"79496525",
x"7937654B",
x"791D656D",
x"7907658E",
x"78FD65B1",
x"790365D8",
x"79186606",
x"793A663B",
x"79636676",
x"798E66B2",
x"79B866F0",
x"79DF672B",
x"7A046760",
x"7A2E678E",
x"7A6367B7",
x"7AAB67D6",
x"7B0D67F2",
x"7B8A6809",
x"7C23681B",
x"7CCE682D",
x"7D83683A",
x"7E316844",
x"7EC66848",
x"7F316848",
x"7F636842",
x"7F526838",
x"7EFA682A",
x"7E5F681A",
x"7D8D6809",
x"7C9467F5",
x"7B8E67DF",
x"7A9367C2",
x"79BB679B",
x"791D6766",
x"78C46720",
x"78B866C5",
x"78F36653",
x"796965D0",
x"7A03653C",
x"7AA764A0",
x"7B3B6403",
x"7BA3636C",
x"7BCE62E2",
x"7BB1626D",
x"7B4C6211",
x"7AAA61CF",
x"79DC61A5",
x"78FC6194",
x"78266198",
x"777361AF",
x"76F661D6",
x"76BE620B",
x"76C9624E",
x"7714629B",
x"778D62F4",
x"78206355",
x"78B463BB",
x"79376423",
x"79966484",
x"79C964DF",
x"79D1652A",
x"79B26565",
x"797D658D",
x"794265A5",
x"791165AE",
x"78F765AE",
x"78F965A5",
x"79116595",
x"7931657F",
x"793F6556",
x"791B6514",
x"78A464AA",
x"77B7640A",
x"763B6325",
x"742461F3",
x"71736072",
x"6E3B5EA9",
x"6AA15CAC",
x"66D85A95",
x"631D5885",
x"5FB056A4",
x"5CCD5515",
x"5AAA53FA",
x"596B5367",
x"59215368",
x"59CF53FA",
x"5B5E550B",
x"5DA95681",
x"6083583A",
x"63BA5A14",
x"67165BEE",
x"6A6C5DAB",
x"6D945F38",
x"7075608A",
x"72FD619D",
x"75286276",
x"76F6631B",
x"78706398",
x"799E63F4",
x"7A8D6439",
x"7B45646D",
x"7BD16493",
x"7C3864AF",
x"7C8064C5",
x"7CB264D6",
x"7CD564E9",
x"7CF06500",
x"7D0D6521",
x"7D2F654F",
x"7D5F658B",
x"7D9E65D6",
x"7DEF6630",
x"7E4C6693",
x"7EB566FC",
x"7F246769",
x"7F9067D6",
x"7FF46844",
x"804F68B1",
x"809B691D",
x"80D9698A",
x"810C69F9",
x"81346A66",
x"81566AD1",
x"81736B32",
x"818D6B86",
x"81A76BC4",
x"81BE6BE8",
x"81D56BEC",
x"81E96BD2",
x"81FE6B9C",
x"82176B4F",
x"82356AF5",
x"825F6A99",
x"82986A42",
x"82E469FD",
x"834869D2",
x"83BC69C2",
x"844169D1",
x"84CB69F9",
x"854F6A34",
x"85C46A77",
x"861D6ABA",
x"86506AF0",
x"865C6B14",
x"86426B20",
x"860A6B11",
x"85C26AED",
x"857B6ABB",
x"85456A86",
x"85326A58",
x"85496A3D",
x"85906A3D",
x"85FD6A59",
x"86836A91",
x"870D6AE1",
x"87816B38",
x"87C86B8D",
x"87CF6BD2",
x"87886BFC",
x"86F76C03",
x"86276BE6",
x"85286BAA",
x"841B6B57",
x"831B6AF9",
x"82436A9C",
x"81AA6A49",
x"81536A09",
x"814169D9",
x"816269B8",
x"81A0699C",
x"81E0697A",
x"82076948",
x"820068FD",
x"81B96897",
x"81346814",
x"8073677D",
x"7F8966DB",
x"7E8A6638",
x"7D9065A3",
x"7CB16525",
x"7C0064C5",
x"7B876487",
x"7B4C646A",
x"7B49646A",
x"7B776484",
x"7BC964B1",
x"7C3464EC",
x"7CA56532",
x"7D176586",
x"7D8065E5",
x"7DDB6652",
x"7E2566CE",
x"7E5F6758",
x"7E8967EC",
x"7E9E6881",
x"7EA1690C",
x"7E89697F",
x"7E5069C8",
x"7DF069D9",
x"7D6069A6",
x"7C996926",
x"7B986858",
x"7A656748",
x"790A6606",
x"779E64AD",
x"7642635A",
x"751D6235",
x"7456615F",
x"741B60F7",
x"748E6117",
x"75CE61C8",
x"77E0630E",
x"7AC564DA",
x"7E636719",
x"829869AA",
x"87356C69",
x"8C046F35",
x"90D871EF",
x"9583747F",
x"99E976D4",
x"9DFA78E8",
x"A1B27ABE",
x"A51B7C5E",
x"A8437DD4",
x"AB407F2B",
x"AE1E8070",
x"B0EB81AC",
x"B3AB82E3",
x"B6578417",
x"B8EA8546",
x"BB538670",
x"BD85878F",
x"BF7588A1",
x"C11B89A4",
x"C2748A93",
x"C3848B6D",
x"C4538C32",
x"C4EB8CE3",
x"C55D8D7B",
x"C5B68E00",
x"C5FF8E70",
x"C6478ECF",
x"C6968F1E",
x"C6F58F66",
x"C7688FAB",
x"C7F88FF3",
x"C8AA9045",
x"C98590A8",
x"CA8C911E",
x"CBC691AD",
x"CD359253",
x"CED79314",
x"D0A993ED",
x"D2A394DE",
x"D4B995E0",
x"D6DA96F3",
x"D8F79810",
x"DAFC9933",
x"DCDC9A54",
x"DE899B6B",
x"DFFB9C6F",
x"E1319D57",
x"E22D9E19",
x"E2F69EB0",
x"E3939F13",
x"E40B9F41",
x"E45E9F38",
x"E48F9EF9",
x"E4959E89",
x"E4679DEE",
x"E3FC9D2E",
x"E34D9C57",
x"E2589B6F",
x"E1299A86",
x"DFCD99A9",
x"DE6298E1",
x"DD09983B",
x"DBE497C1",
x"DB0E9775",
x"DA9C9758",
x"DA959768",
x"DAEF979B",
x"DB9897E9",
x"DC689841",
x"DD3B9897",
x"DDE898DF",
x"DE50990F",
x"DE5A9920",
x"DDFF9911",
x"DD4698E9",
x"DC3E98AA",
x"DB05985C",
x"D9B6980A",
x"D86D97BA",
x"D7409770",
x"D6419733",
x"D5759703",
x"D4DD96E4",
x"D47496D2",
x"D42F96CF",
x"D40596DB",
x"D3EE96F3",
x"D3E29714",
x"D3DE973D",
x"D3DE9768",
x"D3DF978F",
x"D3E197B0",
x"D3E497C5",
x"D3E597D1",
x"D3E797D2",
x"D3E897CE",
x"D3EE97CC",
x"D3F897D5",
x"D40997F0",
x"D4269820",
x"D44A9868",
x"D47698C1",
x"D4A79923",
x"D4D89985",
x"D50399DA",
x"D5259A19",
x"D5399A40",
x"D53D9A4E",
x"D52F9A4B",
x"D50B9A3D",
x"D4C79A2B",
x"D4559A1A",
x"D39D9A02",
x"D27F99D1",
x"D0D79969",
x"CE7798A7",
x"CB3A975E",
x"C7029565",
x"C1C2929D",
x"BB7F8EF9",
x"B45A8A80",
x"AC918552",
x"A4717FAB",
x"9C5D79D6",
x"94BC7429",
x"8DF46EFF",
x"885A6AAA",
x"842E6768",
x"8196655F",
x"8097649B",
x"811B650D",
x"82F7668A",
x"85ED68D9",
x"89BB6BBA",
x"8E1E6EE8",
x"92DC7227",
x"97C5754D",
x"9CB5783A",
x"A1977AE1",
x"A65A7D41",
x"AAF67F64",
x"AF5D815A",
x"B38B8332",
x"B76E84F6",
x"BAF886A9",
x"BE1E884C",
x"C0D189DA",
x"C3128B4B",
x"C4E48C94",
x"C6548DB4",
x"C77C8EA8",
x"C8778F74",
x"C9609024",
x"CA5190C4",
x"CB5E915D",
x"CC9091FD",
x"CDE592AB",
x"CF519366",
x"D0BE942B",
x"D21894F0",
x"D34395A7",
x"D42C9641",
x"D4C696B3",
x"D50596EF",
x"D4EB96EF",
x"D47996B0",
x"D3B99634",
x"D2AD9580",
x"D165949B",
x"CFE89394",
x"CE469277",
x"CC8F9156",
x"CADD9044",
x"C94A8F53",
x"C7FB8E9B",
x"C7138E2C",
x"C6B58E1A",
x"C6F88E6A",
x"C7EB8F1E",
x"C985902D",
x"CBAF917F",
x"CE3992F3",
x"D0E89465",
x"D37995AA",
x"D5AD969D",
x"D74B9720",
x"D82E9723",
x"D84D96AA",
x"D7B095C5",
x"D67B9497",
x"D4E19348",
x"D31C9207",
x"D16790FE",
x"CFF1904F",
x"CEDD900D",
x"CE3A9038",
x"CE0C90C7",
x"CE43919A",
x"CEC69296",
x"CF7F9396",
x"D057947A",
x"D13C952F",
x"D22095AA",
x"D2FF95EA",
x"D3D895FC",
x"D4AA95EF",
x"D56F95D8",
x"D62295C9",
x"D6BC95D5",
x"D7309602",
x"D7799654",
x"D79296C7",
x"D77F9755",
x"D74D97F3",
x"D7099894",
x"D6CD992D",
x"D6AF99B4",
x"D6BE9A20",
x"D70B9A6E",
x"D7929A9A",
x"D84A9AA7",
x"D91F9A99",
x"D9F49A75",
x"DAA49A42",
x"DB129A07",
x"DB1F99C8",
x"DAB69985",
x"D9CB9938",
x"D85F98DA",
x"D67C9858",
x"D43197A1",
x"D19596A3",
x"CEC0954C",
x"CBCA9396",
x"C8C6917F",
x"C5C48F13",
x"C2D08C69",
x"BFF189A5",
x"BD2A86EC",
x"BA7D8466",
x"B7E78236",
x"B5648074",
x"B2EE7F29",
x"B07B7E4F",
x"ADFB7DC7",
x"AB5C7D6D",
x"A87D7D0E",
x"A5457C74",
x"A1947B6B",
x"9D4D79CE",
x"985D7785",
x"92C0748B",
x"8C8170F2",
x"85C26CE1",
x"7EBA688D",
x"77AE6435",
x"70F2601D",
x"6ADF5C82",
x"65C4599A",
x"61E55787",
x"5F69565C",
x"5E615614",
x"5EBD5699",
x"605257C9",
x"62E35975",
x"66235B6E",
x"69C45D83",
x"6D7A5F8D",
x"710C616F",
x"744B6314",
x"7721647A",
x"798765A1",
x"7B876696",
x"7D356768",
x"7EA86828",
x"7FFC68E6",
x"814369B0",
x"82936A8D",
x"83F46B80",
x"85706C87",
x"87036DA0",
x"88A86EBE",
x"8A5A6FD8",
x"8C0D70E5",
x"8DB171D8",
x"8F3B72AB",
x"909E7358",
x"91CF73DF",
x"92C97444",
x"9388748C",
x"941474C6",
x"947474FB",
x"94B5753A",
x"94E7758C",
x"951A75F6",
x"95567679",
x"95A5770D",
x"960A77A6",
x"96807833",
x"970178A2",
x"978878E5",
x"980D78F1",
x"988D78C3",
x"99077861",
x"998477D8",
x"9A0A773D",
x"9AA276A6",
x"9B55762C",
x"9C2575DE",
x"9D1475CD",
x"9E1875FB",
x"9F2B7665",
x"A03C76FE",
x"A14277B4",
x"A2327875",
x"A30A792F",
x"A3CD79D3",
x"A4887A60",
x"A54D7AD8",
x"A6357B4A",
x"A7577BCA",
x"A8CF7C72",
x"AAAE7D5A",
x"AD027E96",
x"AFD38033",
x"B31B8236",
x"B6C98492",
x"BAC48732",
x"BEEA89F3",
x"C3118CAC",
x"C70B8F35",
x"CAAA9165",
x"CDC6931A",
x"D03A9444",
x"D1F494DB",
x"D2E794E6",
x"D31C947D",
x"D2A693BE",
x"D1A492CE",
x"D04091CC",
x"CE9F90DC",
x"CCE8900E",
x"CB3D8F6D",
x"C9AF8EFA",
x"C8468EA7",
x"C6FE8E63",
x"C5CA8E18",
x"C4988DB5",
x"C3538D2A",
x"C1EB8C6D",
x"C05A8B7D",
x"BE9E8A62",
x"BCC28929",
x"BAD887E4",
x"B8FB86A9",
x"B745858B",
x"B5D0849F",
x"B4B883F6",
x"B409839B",
x"B3CE8395",
x"B40783E6",
x"B4A68488",
x"B5998571",
x"B6C78691",
x"B81187D0",
x"B9548914",
x"BA718A43",
x"BB4A8B43",
x"BBC78BFB",
x"BBD68C5A",
x"BB6D8C53",
x"BA878BE3",
x"B9238B0B",
x"B74989D8",
x"B4F88852",
x"B2358688",
x"AEFF8488",
x"AB57825A",
x"A7388007",
x"A2A87D94",
x"9DB17B02",
x"9867785A",
x"92F075A5",
x"8D7A72F4",
x"8842705B",
x"83876DF8",
x"7F8A6BE5",
x"7C836A3E",
x"7A98691D",
x"79DF688D",
x"7A516894",
x"7BD16926",
x"7E2A6A2D",
x"81206B8C",
x"846A6D1A",
x"87C66EB7",
x"8B00703E",
x"8DEF719A",
x"908072BD",
x"92B873AA",
x"94A7746F",
x"966C7520",
x"982B75DB",
x"9A0576BD",
x"9C1A77E1",
x"9E787957",
x"A1287B2A",
x"A4257D56",
x"A7617FC9",
x"AAC58270",
x"AE388527",
x"B19E87C9",
x"B4E08A35",
x"B7E68C46",
x"BA9D8DE7",
x"BCFB8F0A",
x"BEF88FA8",
x"C0938FD1",
x"C1D18F93",
x"C2BD8F11",
x"C3648E6F",
x"C3DA8DD2",
x"C4348D5D",
x"C4888D2E",
x"C4EA8D56",
x"C56A8DDC",
x"C6138EB5",
x"C6ED8FCF",
x"C7F2910D",
x"C91B924B",
x"CA5A9366",
x"CBA0943F",
x"CCDB94C4",
x"CDFE94EA",
x"CEFE94B5",
x"CFDA9437",
x"D093938C",
x"D13392D5",
x"D1C69237",
x"D25891D2",
x"D2F791BC",
x"D3A79207",
x"D46C92B2",
x"D54193B4",
x"D61794F6",
x"D6DE965C",
x"D78397C7",
x"D7F79916",
x"D82E9A2E",
x"D8299AF8",
x"D7EB9B64",
x"D7899B6C",
x"D7189B13",
x"D6B19A5C",
x"D66E9958",
x"D65E9810",
x"D6869697",
x"D6E194FA",
x"D758934B",
x"D7CD9194",
x"D8198FE2",
x"D8188E3F",
x"D7AA8CB6",
x"D6BA8B4F",
x"D5478A0E",
x"D35A88F9",
x"D10E8811",
x"CE888759",
x"CBF486CD",
x"C97B866C",
x"C73D862F",
x"C5508614",
x"C3B98612",
x"C26F8625",
x"C15A8643",
x"C0588666",
x"BF468680",
x"BE01868A",
x"BC6F8676",
x"BA7F8639",
x"B83085CA",
x"B58E8523",
x"B2B08442",
x"AFB98328",
x"ACCD81E3",
x"AA118081",
x"A7A67F19",
x"A5A97DC4",
x"A4267C98",
x"A3247BA8",
x"A2987AFF",
x"A2707AA5",
x"A2907A8C",
x"A2D37AA9",
x"A3177AE0",
x"A3337B12",
x"A3087B26",
x"A2807AFE",
x"A1887A8C",
x"A02179C7",
x"9E5278B6",
x"9C317764",
x"99D575EB",
x"97607464",
x"94EF72E8",
x"9298718F",
x"906D7062",
x"8E716F65",
x"8C9D6E8D",
x"8ADC6DCB",
x"89186D04",
x"87346C26",
x"85176B17",
x"82B769CF",
x"800D684E",
x"7D2D669B",
x"7A3164CF",
x"77446309",
x"74996168",
x"7262600D",
x"70C95F14",
x"6FF35E8D",
x"6FEC5E7E",
x"70B05EE0",
x"72275F9E",
x"742F60A1",
x"769961CC",
x"79306301",
x"7BC9642B",
x"7E42653C",
x"80836630",
x"82846709",
x"844B67D5",
x"85E768A6",
x"876F698D",
x"88F66A9A",
x"8A8D6BD7",
x"8C3E6D44",
x"8E076ED9",
x"8FDD708A",
x"91AE723E",
x"936373DC",
x"94E7754E",
x"9627767C",
x"9717775A",
x"97B577DB",
x"980A7806",
x"982877E5",
x"9824778B",
x"981B770D",
x"9829768C",
x"98667622",
x"98E675E5",
x"99B275EA",
x"9AD2763C",
x"9C3D76DE",
x"9DED77CD",
x"9FD378FC",
x"A1DD7A5E",
x"A3FE7BDE",
x"A6237D6A",
x"A8427EF1",
x"AA4C8067",
x"AC3C81C3",
x"AE088300",
x"AFAB8419",
x"B11C850F",
x"B25685E2",
x"B354868D",
x"B40F870E",
x"B4888760",
x"B4BD8780",
x"B4B58767",
x"B47A8718",
x"B4178695",
x"B39E85EA",
x"B3218522",
x"B2B28452",
x"B263838B",
x"B23F82E3",
x"B2538268",
x"B2A68229",
x"B3388226",
x"B4088261",
x"B50F82D1",
x"B643836B",
x"B7968422",
x"B8FA84E7",
x"BA5A85B2",
x"BBA6867B",
x"BCC9873F",
x"BDB287FA",
x"BE5488B1",
x"BEA8895F",
x"BEA68A05",
x"BE548A9D",
x"BDBC8B1F",
x"BCEA8B84",
x"BBF38BC2",
x"BAED8BD3",
x"B9EE8BB5",
x"B90B8B6D",
x"B8538B04",
x"B7D48A88",
x"B7948A0D",
x"B792899E",
x"B7CC894A",
x"B8358915",
x"B8C08900",
x"B95A88FD",
x"B9F188FB",
x"BA6E88E9",
x"BABF88AF",
x"BAD18840",
x"BA9B8794",
x"BA1386AC",
x"B9438597",
x"B835846D",
x"B701834A",
x"B5C3824F",
x"B4A28199",
x"B3BF813F",
x"B336814A",
x"B31E81BB",
x"B37A827E",
x"B4408377",
x"B5568484",
x"B694857B",
x"B7CA863B",
x"B8CD86A7",
x"B97486AF",
x"B9A58659",
x"B95A85AF",
x"B89B84D0",
x"B78183DD",
x"B62E82FA",
x"B4C28240",
x"B35681BF",
x"B1F08175",
x"B084814F",
x"AEEE8126",
x"ACFE80CA",
x"AA738008",
x"A7157EB2",
x"A2BD7CA3",
x"9D5F79D4",
x"970A764D",
x"8FFA7233",
x"88866DBF",
x"8120693B",
x"7A3F64F2",
x"745C612E",
x"6FD45E2C",
x"6CE65C17",
x"6BAB5AFE",
x"6C115AE1",
x"6DDE5BA6",
x"70BE5D27",
x"744C5F31",
x"78216190",
x"7BE06413",
x"7F41668E",
x"821368E1",
x"84446AF2",
x"85D66CB1",
x"86E56E19",
x"87926F2A",
x"88076FE8",
x"8867705C",
x"88CF7094",
x"895270A1",
x"89F67090",
x"8AB87075",
x"8B93705B",
x"8C79704F",
x"8D5F705A",
x"8E3B707C",
x"8F0670B1",
x"8FB870F0",
x"904F712E",
x"90C6715C",
x"9117716F",
x"9139715B",
x"9127711F",
x"90D670B9",
x"90417030",
x"8F666F8F",
x"8E496EE1",
x"8CF36E33",
x"8B716D90",
x"89DC6CFF",
x"88496C83",
x"86D36C1D",
x"85906BCE",
x"84946B92",
x"83EC6B66",
x"839B6B4C",
x"83A16B42",
x"83F66B4F",
x"848E6B75",
x"855D6BB7",
x"86566C19",
x"876D6C9A",
x"889D6D3A",
x"89DF6DF0",
x"8B326EB4",
x"8C916F79",
x"8DFC7037",
x"8F6970E1",
x"90D0716F",
x"922471DC",
x"93527226",
x"9449724D",
x"94F77255",
x"954B7243",
x"953B721A",
x"94C271E1",
x"93E67197",
x"92AE7143",
x"913170E4",
x"8F83707C",
x"8DC37010",
x"8C0D6FA6",
x"8A806F43",
x"89346EEF",
x"883F6EB4",
x"87AF6E96",
x"878D6E9A",
x"87D66EC1",
x"88866F08",
x"898A6F64",
x"8AD06FCB",
x"8C3F7033",
x"8DBF708F",
x"8F3570D2",
x"908A70FB",
x"91A77105",
x"927E70F4",
x"930470CD",
x"93367099",
x"9314705F",
x"92A77026",
x"91FA6FEF",
x"911D6FBB",
x"90216F88",
x"8F1A6F4D",
x"8E1B6F06",
x"8D386EB3",
x"8C7D6E52",
x"8BF96DEC",
x"8BAF6D8A",
x"8BA26D37",
x"8BCE6D00",
x"8C276CF0",
x"8C9E6D0D",
x"8D256D57",
x"8DA86DC5",
x"8E186E4E",
x"8E696EDF",
x"8E946F69",
x"8E9A6FDC",
x"8E7D7030",
x"8E48705F",
x"8E017069",
x"8DB17055",
x"8D577029",
x"8CEF6FE8",
x"8C676F94",
x"8BAA6F26",
x"8A9E6E90",
x"89286DC7",
x"87326CB5",
x"84AF6B51",
x"81A26991",
x"7E1E677F",
x"7A42652A",
x"764162AF",
x"72516039",
x"6EAD5DF0",
x"6B8A5C00",
x"69195A8B",
x"677559A9",
x"66AB5963",
x"66BB59AE",
x"678D5A76",
x"69055B9A",
x"6AFA5CF4",
x"6D455E62",
x"6FBC5FC3",
x"723E6103",
x"74AE6217",
x"76F96303",
x"791163D0",
x"7AF36491",
x"7C9E6558",
x"7E1B6634",
x"7F726732",
x"80B16858",
x"81E569A1",
x"831E6B07",
x"84676C7C",
x"85CE6DEF",
x"87556F52",
x"88FC7096",
x"8ABE71B4",
x"8C8D72A4",
x"8E597366",
x"901073FE",
x"919A746B",
x"92E674B4",
x"93E674DB",
x"949274E4",
x"94EC74CE",
x"94F97499",
x"94C67448",
x"946973DC",
x"93F4735A",
x"937B72C8",
x"93147233",
x"92C971A4",
x"92A4712B",
x"92AA70D8",
x"92D970B4",
x"932C70C5",
x"939E7113",
x"94257196",
x"94BB7247",
x"955A7319",
x"960073FC",
x"96AC74E0",
x"976075B4",
x"9821766F",
x"98F1770B",
x"99D97783",
x"9AD977E0",
x"9BEE7829",
x"9D177867",
x"9E4878A6",
x"9F7678EE",
x"A08E7943",
x"A18179A5",
x"A23F7A0F",
x"A2BD7A77",
x"A2F77AD4",
x"A2ED7B1F",
x"A2AE7B4E",
x"A24A7B61",
x"A1DF7B5B",
x"A1837B41",
x"A1527B20",
x"A1617B02",
x"A1B97AF2",
x"A25A7AF9",
x"A3397B19",
x"A43B7B51",
x"A5427B9B",
x"A6297BED",
x"A6D27C3A",
x"A71C7C75",
x"A6F87C96",
x"A65E7C92",
x"A5537C64",
x"A3E67C09",
x"A22C7B85",
x"A0457ADA",
x"9E467A09",
x"9C4B791B",
x"9A607815",
x"989376FE",
x"96E375E1",
x"955274C8",
x"93DC73C0",
x"927D72D7",
x"91347219",
x"9001718F",
x"8EED713D",
x"8DFD7120",
x"8D397133",
x"8CAB7162",
x"8C507199",
x"8C2B71C1",
x"8C2E71C4",
x"8C4F718F",
x"8C797117",
x"8C9B705C",
x"8CA56F66",
x"8C8A6E4B",
x"8C436D23",
x"8BD36C09",
x"8B3F6B19",
x"8A956A68",
x"89E36A04",
x"893869ED",
x"889B6A1C",
x"88136A7A",
x"879A6AEC",
x"87276B52",
x"86A86B8D",
x"860B6B83",
x"853A6B23",
x"84246A65",
x"82BF694E",
x"810A67ED",
x"7F0D6660",
x"7CDA64C4",
x"7A8D633B",
x"784261E6",
x"761B60E0",
x"7435603C",
x"72AB6003",
x"718E602F",
x"70E960B7",
x"70BB6183",
x"71016277",
x"71AE637C",
x"72B46473",
x"7400654B",
x"758665F5",
x"77386670",
x"790D66C2",
x"7AFE66FC",
x"7D096731",
x"7F2A6779",
x"816067E9",
x"83AF6894",
x"86116980",
x"88866AB0",
x"8B066C16",
x"8D886DA4",
x"90046F3E",
x"926F70CE",
x"94B97239",
x"96DA736C",
x"98C5745B",
x"9A6D7505",
x"9BCF7571",
x"9CE675AD",
x"9DB375D2",
x"9E3D75F6",
x"9E8B7630",
x"9EAE7690",
x"9EB27722",
x"9EAB77E2",
x"9EA778CB",
x"9EB579CB",
x"9EE07AD0",
x"9F2E7BC1",
x"9F9F7C8B",
x"A0327D20",
x"A0DF7D78",
x"A19F7D95",
x"A26D7D7F",
x"A3407D49",
x"A4177D04",
x"A4EE7CC4",
x"A5C87C9E",
x"A6A87C9C",
x"A7927CC9",
x"A88B7D1F",
x"A9917D98",
x"AAA37E26",
x"ABBC7EB7",
x"ACD27F36",
x"ADD67F98",
x"AEBD7FCD",
x"AF787FCF",
x"AFFB7FA0",
x"B03C7F47",
x"B0367ED3",
x"AFEB7E50",
x"AF637DD3",
x"AEA97D6D",
x"ADCC7D2C",
x"ACE17D1C",
x"ABF87D3F",
x"AB257D91",
x"AA787E07",
x"A9FD7E94",
x"A9BB7F23",
x"A9B67FA5",
x"A9ED8005",
x"AA5C8039",
x"AAFB8039",
x"ABC58007",
x"ACAC7FA9",
x"ADA87F32",
x"AEB27EB6",
x"AFC07E47",
x"B0C97DFB",
x"B1C57DE1",
x"B2AD7E01",
x"B37D7E5B",
x"B42D7EE7",
x"B4BF7F91",
x"B52F8046",
x"B57B80EE",
x"B5A58170",
x"B5AB81B7",
x"B58781B7",
x"B533816A",
x"B4A580CF",
x"B3D27FF0",
x"B2A97EDB",
x"B1237DA0",
x"AF3C7C56",
x"ACF47B0C",
x"AA5979D4",
x"A77F78B7",
x"A48B77BE",
x"A1A276EE",
x"9EEE7646",
x"9C9575C1",
x"9AB4755A",
x"99577506",
x"987E74C0",
x"98137479",
x"97F47429",
x"97F973C8",
x"97F37350",
x"97BB72BE",
x"97337213",
x"96527155",
x"9518708C",
x"939C6FC4",
x"91FA6F09",
x"90526E68",
x"8EC36DE8",
x"8D5F6D8A",
x"8C286D4D",
x"8B0E6D21",
x"89F36CF9",
x"88AE6CBA",
x"87126C4A",
x"84FB6B94",
x"82506A86",
x"7F116919",
x"7B526751",
x"773F653E",
x"73186301",
x"6F2860C2",
x"6BBB5EAC",
x"69165CED",
x"67695BA9",
x"66CF5AFD",
x"674A5AF1",
x"68BD5B81",
x"6AF65C95",
x"6DB75E08",
x"70B25FAE",
x"73A76153",
x"765562CE",
x"789163FA",
x"7A4264C2",
x"7B696525",
x"7C13652F",
x"7C6364FD",
x"7C8364B2",
x"7CA16479",
x"7CE56476",
x"7D7064C8",
x"7E55657D",
x"7F966697",
x"81256806",
x"82EC69AA",
x"84C66B5F",
x"868E6CFA",
x"88246E55",
x"896D6F54",
x"8A5C6FE2",
x"8AF17002",
x"8B3B6FBE",
x"8B536F34",
x"8B5A6E89",
x"8B736DE5",
x"8BBB6D6E",
x"8C496D42",
x"8D276D78",
x"8E4F6E12",
x"8FB76F0A",
x"9143704A",
x"92DA71B4",
x"94607327",
x"95BE7483",
x"96E775AD",
x"97D87690",
x"98977729",
x"99357779",
x"99C6778F",
x"9A64777E",
x"9B24775B",
x"9C15773E",
x"9D427737",
x"9EA87755",
x"A0407799",
x"A1FB7802",
x"A3C57888",
x"A584791D",
x"A72679B7",
x"A8947A47",
x"A9C07AC4",
x"AA9C7B29",
x"AB237B71",
x"AB537B9C",
x"AB2F7BAD",
x"AABF7BA9",
x"AA0B7B93",
x"A9257B6E",
x"A8197B40",
x"A6FF7B0C",
x"A5EA7ADA",
x"A4ED7AAC",
x"A41B7A8C",
x"A3857A7E",
x"A3387A86",
x"A3387AA8",
x"A3857AE0",
x"A41A7B2A",
x"A4E77B7E",
x"A5DD7BD0",
x"A6E77C13",
x"A7F37C3C",
x"A8EB7C44",
x"A9C67C28",
x"AA767BE8",
x"AAF87B8C",
x"AB4C7B22",
x"AB717AB3",
x"AB6A7A50",
x"AB3879FE",
x"AAD779C4",
x"AA47799F",
x"A9827988",
x"A8817971",
x"A742794D",
x"A5C3790E",
x"A40B78A7",
x"A2257816",
x"A0227758",
x"9E157675",
x"9C177579",
x"9A3B7472",
x"9895736F",
x"972F727E",
x"961071A7",
x"953270EE",
x"948D7052",
x"940E6FCF",
x"93A76F5C",
x"93456EF0",
x"92DA6E86",
x"925F6E19",
x"91CE6DAB",
x"912C6D41",
x"90836CE2",
x"8FD96C97",
x"8F396C66",
x"8EAA6C57",
x"8E2C6C63",
x"8DBC6C86",
x"8D4B6CAE",
x"8CC26CC7",
x"8C096CBA",
x"8B036C6F",
x"89956BD2",
x"87AA6AD7",
x"85356977",
x"823967BB",
x"7EC665B4",
x"7AFA6379",
x"7704612B",
x"731A5EEE",
x"6F775CE3",
x"6C585B26",
x"69ED59D3",
x"685C58F3",
x"67BB588C",
x"6807589B",
x"692E5912",
x"6B0C59E3",
x"6D705AF8",
x"70275C3F",
x"72FC5DA4",
x"75C25F18",
x"785B608D",
x"7AAF61FA",
x"7CBC6359",
x"7E8A64A4",
x"802865DB",
x"81AE66FA",
x"832F6804",
x"84C268F9",
x"867169D9",
x"88426AA7",
x"8A376B66",
x"8C466C1A",
x"8E696CC8",
x"90936D73",
x"92B66E20",
x"94CC6ED4",
x"96CB6F92",
x"98A8705B",
x"9A617130",
x"9BED7210",
x"9D4972F9",
x"9E6E73EB",
x"9F5A74E1",
x"A00F75DB",
x"A09276D7",
x"A0ED77D2",
x"A12F78D1",
x"A16A79CE",
x"A1B57ACB",
x"A2257BC4",
x"A2CF7CB4",
x"A3BD7D98",
x"A4F77E67",
x"A6777F16",
x"A82E7FA5",
x"AA05800A",
x"ABE38045",
x"ADA68054",
x"AF388043",
x"B07D8019",
x"B16B7FE6",
x"B1FE7FB7",
x"B23D7F9F",
x"B2377FAC",
x"B2057FE6",
x"B1C28050",
x"B18580EB",
x"B16781AD",
x"B177828A",
x"B1BD836E",
x"B23B8449",
x"B2EA8507",
x"B3C0859E",
x"B4B28604",
x"B5B88638",
x"B6CA863F",
x"B7E78623",
x"B91285F7",
x"BA4E85C9",
x"BBA385AC",
x"BD1285B1",
x"BE9985DD",
x"C032863B",
x"C1CA86C6",
x"C34E877A",
x"C4A3884A",
x"C5B2892B",
x"C6608A0A",
x"C69C8ADA",
x"C6638B8E",
x"C5B38C1D",
x"C49F8C7E",
x"C33D8CAF",
x"C1AB8CAE",
x"C0088C7D",
x"BE778C1E",
x"BD0E8B97",
x"BBE38AEC",
x"BAFB8A22",
x"BA548942",
x"B9E68852",
x"B99E8759",
x"B9668660",
x"B92C8571",
x"B8DE8492",
x"B87283CF",
x"B7E68329",
x"B73882A6",
x"B6738247",
x"B59E8208",
x"B4C481E1",
x"B3EB81C9",
x"B31281B3",
x"B230818F",
x"B13D8153",
x"B02880F2",
x"AEE38067",
x"AD667FAF",
x"ABAC7ECF",
x"A9BC7DCD",
x"A7A57CB7",
x"A5807B9C",
x"A3647A89",
x"A1707989",
x"9FB378A3",
x"9E3977D5",
x"9CFB771D",
x"9BEA766E",
x"9AE675BA",
x"99CA74F1",
x"98747408",
x"96C372F5",
x"94A771B7",
x"921B7052",
x"8F316ED7",
x"8C066D54",
x"88C66BE1",
x"85A76A94",
x"82D86980",
x"808668B4",
x"7ED3683A",
x"7DD36810",
x"7D8D6835",
x"7DF6689D",
x"7EFF693F",
x"80936A0D",
x"82986AFF",
x"84FD6C0D",
x"87B26D35",
x"8AAA6E79",
x"8DDF6FD8",
x"914B715A",
x"94E972FC",
x"98AC74C1",
x"9C8A76A5",
x"A06B789F",
x"A4397AA2",
x"A7D67CA0",
x"AB257E8C",
x"AE098056",
x"B07781F4",
x"B2618363",
x"B3CE84A2",
x"B4CE85B9",
x"B57D86B8",
x"B5FA87AC",
x"B66B88A9",
x"B6F389BE",
x"B7A88AF3",
x"B8988C49",
x"B9C08DB8",
x"BB128F2F",
x"BC719096",
x"BDC091CF",
x"BEDD92BF",
x"BFAF934F",
x"C0289373",
x"C04A9327",
x"C0269279",
x"BFDB917F",
x"BF919059",
x"BF6B8F2F",
x"BF8C8E24",
x"C00E8D56",
x"C0F28CDD",
x"C2368CC1",
x"C3C08D01",
x"C56E8D93",
x"C71F8E62",
x"C8AD8F58",
x"C9FF905C",
x"CB02915D",
x"CBAF9249",
x"CC099317",
x"CC1993C1",
x"CBEB9441",
x"CB889496",
x"CAF794BF",
x"CA3694BA",
x"C9479482",
x"C8239417",
x"C6CB937D",
x"C54792B9",
x"C3A291D8",
x"C1F490E7",
x"C05B9000",
x"BEFE8F35",
x"BDFC8E9D",
x"BD748E48",
x"BD7A8E41",
x"BE118E86",
x"BF2D8F13",
x"C0B78FD6",
x"C28890BB",
x"C47191AB",
x"C640928D",
x"C7C7934B",
x"C8E093D5",
x"C96B9420",
x"C9589425",
x"C8A693E3",
x"C758935B",
x"C5849291",
x"C340918D",
x"C0AC9053",
x"BDE78EED",
x"BB118D66",
x"B84A8BC6",
x"B5AB8A1E",
x"B349887A",
x"B13386E9",
x"AF738578",
x"AE058433",
x"ACE6831F",
x"AC05823D",
x"AB528185",
x"AAB580F0",
x"AA1E806E",
x"A97A7FF2",
x"A8BC7F6E",
x"A7DF7ED9",
x"A6E07E2C",
x"A5C67D6A",
x"A49C7C99",
x"A36E7BC4",
x"A24A7AF9",
x"A13F7A47",
x"A05979B7",
x"9FA27958",
x"9F24792C",
x"9EE77936",
x"9EEE7974",
x"9F3879DE",
x"9FBC7A68",
x"A06A7B01",
x"A1227B92",
x"A1BE7BFF",
x"A2047C29",
x"A1B87BEE",
x"A0977B2C",
x"9E6779C4",
x"9AFB77A5",
x"964274C7",
x"90487135",
x"893C6D0F",
x"81736886",
x"795F63DD",
x"71845F5F",
x"6A6C5B5C",
x"64995818",
x"607355CF",
x"5E3F549F",
x"5E1A5494",
x"5FF35599",
x"63925788",
x"689E5A26",
x"6EB05D35",
x"75586076",
x"7C2D63B2",
x"82D666C8",
x"8915699E",
x"8EBE6C33",
x"93BC6E8C",
x"980F70BA",
x"9BC372CB",
x"9EE374C8",
x"A18376B4",
x"A3AF7888",
x"A5717A33",
x"A6D27BA5",
x"A7D37CCA",
x"A87D7D96",
x"A8D47E08",
x"A8E67E28",
x"A8BD7E07",
x"A8697DBF",
x"A7F77D6A",
x"A7777D20",
x"A6F37CF7",
x"A6717CF1",
x"A5F67D0F",
x"A5817D41",
x"A5117D78",
x"A4A57D9B",
x"A43B7D99",
x"A3D37D64",
x"A36D7CFC",
x"A30C7C65",
x"A2B27BAF",
x"A2607AEF",
x"A21C7A3E",
x"A1E679B0",
x"A1BE7957",
x"A1A67939",
x"A1A17958",
x"A1AC79AD",
x"A1C97A2A",
x"A1F47AC0",
x"A22C7B5E",
x"A26E7BF8",
x"A2B67C84",
x"A2FE7CFF",
x"A33D7D6A",
x"A3717DC7",
x"A3927E1C",
x"A39C7E70",
x"A38B7EC0",
x"A35D7F0A",
x"A3127F49",
x"A2A67F72",
x"A21B7F77",
x"A16B7F4D",
x"A09B7EEB",
x"9FA77E4A",
x"9E957D6F",
x"9D6A7C65",
x"9C337B3A",
x"9B047A06",
x"99ED78E2",
x"990A77E5",
x"98717725",
x"983B76AF",
x"9874768B",
x"992876B7",
x"9A56772A",
x"9BF477D8",
x"9DF378AF",
x"A03B799D",
x"A2B37A95",
x"A5427B8B",
x"A7CF7C7C",
x"AA437D65",
x"AC8F7E49",
x"AE9F7F25",
x"B06A7FFC",
x"B1E480C9",
x"B3028184",
x"B3BD8223",
x"B411829C",
x"B40182E4",
x"B39282F6",
x"B2D682D0",
x"B1DE827B",
x"B0CC8205",
x"AFBA8182",
x"AECC8108",
x"AE1E80AF",
x"ADC68087",
x"ADD3809C",
x"AE4A80F5",
x"AF28818E",
x"B059825D",
x"B1CC8350",
x"B3668459",
x"B50B8563",
x"B6A28662",
x"B8168748",
x"B9578812",
x"BA5D88C0",
x"BB258956",
x"BBB989DC",
x"BC288A5A",
x"BC888ADC",
x"BCF18B69",
x"BD788C06",
x"BE2D8CB2",
x"BF128D67",
x"C0188E1A",
x"C11B8EB1",
x"C1E78F13",
x"C2378F1D",
x"C1BF8EAB",
x"C0308D9B",
x"BD4D8BD3",
x"B8EE8942",
x"B30C85E6",
x"ABCA81D1",
x"A36D7D2C",
x"9A5D7826",
x"911F7305",
x"883C6E12",
x"803C6996",
x"799065D0",
x"748962F0",
x"71516111",
x"6FE36038",
x"70196050",
x"71A46134",
x"742A62AB",
x"773F647A",
x"7A836665",
x"7DA16831",
x"805969B8",
x"82866ADC",
x"841B6B96",
x"85256BEB",
x"85BE6BEC",
x"860A6BB7",
x"86346B6B",
x"86636B27",
x"86B76B06",
x"87466B19",
x"881B6B65",
x"89326BEB",
x"8A816C9C",
x"8BF36D66",
x"8D6D6E35",
x"8ED76EF5",
x"901A6F90",
x"91226FFF",
x"91E4703B",
x"925A7047",
x"928B702B",
x"927E6FF5",
x"92406FB0",
x"91E06F68",
x"916A6F24",
x"90E36EE9",
x"90506EB5",
x"8FAC6E83",
x"8EF36E4D",
x"8E1A6E0D",
x"8D1D6DBF",
x"8BF76D66",
x"8AAF6D04",
x"894F6CA6",
x"87E96C52",
x"86906C16",
x"855C6BF9",
x"84656C02",
x"83B86C2D",
x"835F6C78",
x"83566CD7",
x"83956D3E",
x"840D6D9E",
x"84A76DEF",
x"85506E24",
x"85F66E3D",
x"868E6E38",
x"87146E20",
x"87906DFA",
x"880A6DD9",
x"88946DC5",
x"893E6DCB",
x"8A136DF3",
x"8B176E3F",
x"8C486EB0",
x"8D956F3B",
x"8EE96FD4",
x"9024706B",
x"912570EC",
x"91D07147",
x"920D716B",
x"91D0714E",
x"911770E9",
x"8FF27044",
x"8E796F65",
x"8CD06E62",
x"8B1F6D4E",
x"898E6C42",
x"883F6B57",
x"874B6A9D",
x"86C16A26",
x"86A169F2",
x"86E06A03",
x"87676A4B",
x"881E6ABD",
x"88E66B47",
x"89A76BD5",
x"8A4B6C5B",
x"8AC96CCD",
x"8B1F6D28",
x"8B586D6E",
x"8B7F6DA4",
x"8BA76DD7",
x"8BE06E0D",
x"8C396E57",
x"8CBC6EB7",
x"8D666F35",
x"8E326FD1",
x"8F147085",
x"8FF67147",
x"90C8720D",
x"917672CA",
x"91F1736C",
x"922F73E6",
x"922E742D",
x"91EF7437",
x"917B73FF",
x"90DD7389",
x"902472DC",
x"8F5D7203",
x"8E95710F",
x"8DD57012",
x"8D216F1C",
x"8C776E3D",
x"8BD26D7C",
x"8B246CD9",
x"8A5A6C4F",
x"89636BD2",
x"88286B4C",
x"869A6AAE",
x"84AB69E5",
x"825C68E6",
x"7FB867B1",
x"7CD6664C",
x"79DF64CC",
x"7701634C",
x"747661EF",
x"727960D5",
x"713B601E",
x"70E95FE0",
x"71986027",
x"734B60F2",
x"75F06234",
x"795F63D8",
x"7D5F65BF",
x"81AE67CF",
x"860969E8",
x"8A2F6BF3",
x"8DF46DDE",
x"91356F9F",
x"93E97134",
x"961872A1",
x"97DD73EE",
x"995C7523",
x"9AC3764B",
x"9C3C7772",
x"9DED789D",
x"9FEE79D7",
x"A2507B26",
x"A5127C8C",
x"A8287E0F",
x"AB7D7FAC",
x"AEF48164",
x"B2748332",
x"B5DE850A",
x"B91E86E0",
x"BC1B88A7",
x"BECB8A4D",
x"C1238BC9",
x"C31F8D0D",
x"C4BF8E10",
x"C6018ED1",
x"C6E88F4F",
x"C77A8F90",
x"C7B98F9B",
x"C7AD8F77",
x"C7618F2C",
x"C6E18EC5",
x"C6398E43",
x"C5788DAF",
x"C4AC8D0B",
x"C3E08C5A",
x"C31B8BA1",
x"C25D8AE2",
x"C1A08A1D",
x"C0DD8956",
x"C002888B",
x"BF0287BE",
x"BDD486EA",
x"BC73860F",
x"BAE3852F",
x"B935844A",
x"B7848367",
x"B5F0828C",
x"B49B81C7",
x"B3A38121",
x"B31F80A3",
x"B3128054",
x"B3778033",
x"B42F803C",
x"B5168063",
x"B5FD8099",
x"B6B380CF",
x"B71280F5",
x"B7048105",
x"B68180FD",
x"B59B80E4",
x"B47780CA",
x"B34680C5",
x"B24080E8",
x"B199814D",
x"B17B81FE",
x"B1FB8300",
x"B318844A",
x"B4B985CA",
x"B6B08762",
x"B8C588EC",
x"BAB68A45",
x"BC4E8B4B",
x"BD618BE0",
x"BDDA8BFA",
x"BDBD8B97",
x"BD228AC2",
x"BC388995",
x"BB308831",
x"BA4486BC",
x"B99F855A",
x"B95E842B",
x"B9858346",
x"BA0282B5",
x"BAB2827A",
x"BB63828A",
x"BBE382D0",
x"BC058338",
x"BBAF83A8",
x"BADA840F",
x"B99B8460",
x"B8198494",
x"B68C84AD",
x"B52F84B5",
x"B43884B3",
x"B3CC84B5",
x"B3FA84BD",
x"B4B284CF",
x"B5CC84E1",
x"B70C84EC",
x"B82C84DA",
x"B8E6849E",
x"B901842C",
x"B85A837D",
x"B6EA8291",
x"B4C68172",
x"B2198033",
x"AF247EEA",
x"AC267DA8",
x"A95B7C81",
x"A6F17B7E",
x"A4FA7A9D",
x"A37079D4",
x"A2357910",
x"A1177834",
x"9FD77729",
x"9E3D75D7",
x"9C1A7430",
x"994F7233",
x"95DA6FEB",
x"91D36D73",
x"8D6A6AEF",
x"88DF6889",
x"847C666A",
x"808964BC",
x"7D44639A",
x"7ADB6314",
x"7968632B",
x"78EB63D5",
x"795364F7",
x"7A836673",
x"7C4E6826",
x"7E8969ED",
x"810D6BAD",
x"83B96D4F",
x"867C6ECD",
x"89487023",
x"8C1A715A",
x"8EF6727F",
x"91DD73A3",
x"94D274D5",
x"97CF761F",
x"9ACC7786",
x"9DB97908",
x"A0857A9B",
x"A31E7C30",
x"A5737DB7",
x"A77A7F1C",
x"A9328053",
x"AA9F814F",
x"ABCC820B",
x"ACCC828A",
x"ADAC82D4",
x"AE8182F7",
x"AF578304",
x"B033830C",
x"B116831F",
x"B1FA8346",
x"B2D4838A",
x"B39983EA",
x"B43C8463",
x"B4B584E8",
x"B4FD8571",
x"B51885EE",
x"B50C8653",
x"B4E18698",
x"B4A286B3",
x"B45A86A5",
x"B40F866D",
x"B3C6860F",
x"B37D8595",
x"B32F8504",
x"B2D68463",
x"B26883B9",
x"B1E1830B",
x"B13F825E",
x"B08081B3",
x"AFAB810B",
x"AEC9806A",
x"ADE97FCF",
x"AD147F3C",
x"AC5E7EB7",
x"ABD27E44",
x"AB7D7DEA",
x"AB677DAD",
x"AB9B7D96",
x"AC187DA9",
x"ACDE7DE7",
x"ADE97E50",
x"AF2F7EE0",
x"B0A17F8F",
x"B22D8054",
x"B3BF8126",
x"B54481FA",
x"B6AA82C6",
x"B7E78388",
x"B8F5843C",
x"B9D784E7",
x"BA978591",
x"BB44863F",
x"BBF586FB",
x"BCBA87CF",
x"BDA688B9",
x"BEC189BE",
x"C0128AD5",
x"C1928BFA",
x"C3368D25",
x"C4EE8E4C",
x"C6A68F6A",
x"C84C907D",
x"C9C99180",
x"CB109277",
x"CC13935F",
x"CCC99438",
x"CD2A94FD",
x"CD3395A5",
x"CCE79621",
x"CC479665",
x"CB619660",
x"CA44960A",
x"C907955F",
x"C7C09465",
x"C6899328",
x"C57E91C1",
x"C4AA9045",
x"C41B8ED2",
x"C3C68D7E",
x"C3A08C5C",
x"C38E8B70",
x"C3728ABB",
x"C32D8A34",
x"C2A989CC",
x"C1D88976",
x"C0BD8921",
x"BF6A88C8",
x"BDF58866",
x"BC8287FE",
x"BB2D8792",
x"BA08872B",
x"B91286C2",
x"B8338656",
x"B74385D4",
x"B607852B",
x"B438843D",
x"B19882F2",
x"ADF88137",
x"A9427EFF",
x"A37D7C4E",
x"9CD97932",
x"95A975CD",
x"8E59724B",
x"875F6EDE",
x"81356BBA",
x"7C44690E",
x"78D96701",
x"771D65AA",
x"7710650D",
x"788D6524",
x"7B4E65D8",
x"7EF56709",
x"83236893",
x"87766A52",
x"8BA16C28",
x"8F6E6DFC",
x"92C26FBE",
x"9598716B",
x"98057302",
x"9A2B748C",
x"9C2B760F",
x"9E27778F",
x"A0327910",
x"A2537A8C",
x"A47D7BF7",
x"A6987D43",
x"A8887E60",
x"AA2B7F3C",
x"AB677FD1",
x"AC33801C",
x"AC918022",
x"AC977FF0",
x"AC647F9E",
x"AC287F42",
x"AC127EFA",
x"AC507ED9",
x"AD057EF1",
x"AE447F4A",
x"B0117FE8",
x"B25C80C2",
x"B50281C5",
x"B7D982E0",
x"BAAC83FD",
x"BD4A850A",
x"BF8685F6",
x"C13C86B5",
x"C2578742",
x"C2D6879D",
x"C2C087C8",
x"C22F87CC",
x"C14687B2",
x"C02D8784",
x"BF0F8749",
x"BE14870B",
x"BD5986D2",
x"BCF7869F",
x"BCFA867A",
x"BD5D8660",
x"BE148652",
x"BF02864C",
x"C0088649",
x"C0FB8643",
x"C1B58636",
x"C20F861C",
x"C1EE85F3",
x"C13F85B8",
x"BFFE856D",
x"BE368517",
x"BBFF84BD",
x"B981846A",
x"B6E78425",
x"B46483F8",
x"B22583E7",
x"B05183F6",
x"AF058422",
x"AE528464",
x"AE3384B5",
x"AE9C8508",
x"AF758553",
x"B09E8588",
x"B1F185A2",
x"B34C8598",
x"B491856C",
x"B5A6851B",
x"B67D84AC",
x"B70A8425",
x"B746838A",
x"B73382E1",
x"B6D18230",
x"B61F8178",
x"B51F80BC",
x"B3CE7FFB",
x"B2307F33",
x"B0497E64",
x"AE1B7D89",
x"ABB57CA2",
x"A9227BAC",
x"A6777AA9",
x"A3CC799C",
x"A1347889",
x"9EC67774",
x"9C947667",
x"9AAB756A",
x"990D7485",
x"97BB73C4",
x"96AC732F",
x"95D272C8",
x"951C7293",
x"947A7289",
x"93DA72A3",
x"932E72D4",
x"926C730C",
x"9191733E",
x"909E735C",
x"8F9A735B",
x"8E907337",
x"8D8872EF",
x"8C937288",
x"8BB57208",
x"8AF67179",
x"8A5270E2",
x"89BF7044",
x"892B6F9D",
x"887C6EE6",
x"87946E12",
x"86536D0F",
x"849B6BCE",
x"82556A42",
x"7F736860",
x"7BF4662B",
x"77E663AB",
x"736660F2",
x"6E9D5E1A",
x"69BE5B43",
x"6503588F",
x"60A3561F",
x"5CD1540E",
x"59B7526E",
x"576F514C",
x"560850A6",
x"55795078",
x"55B350B0",
x"5693513F",
x"57F5520B",
x"59AB5304",
x"5B905416",
x"5D7B5533",
x"5F515650",
x"60FF5766",
x"627D586D",
x"63CC5960",
x"64F25A3D",
x"65F95B00",
x"66EF5BA1",
x"67D95C1F",
x"68C15C78",
x"69A65CAB",
x"6A845CBD",
x"6B555CB6",
x"6C115C9F",
x"6CB05C86",
x"6D2D5C76",
x"6D865C7B",
x"6DBF5C9F",
x"6DDF5CE4",
x"6DE95D4B",
x"6DE95DCB",
x"6DE25E59",
x"6DD85EE9",
x"6DCB5F69",
x"6DBA5FCB",
x"6DA16003",
x"6D7A600A",
x"6D475FDD",
x"6D035F81",
x"6CB75EFA",
x"6C685E57",
x"6C1D5DA5",
x"6BDF5CF3",
x"6BB55C52",
x"6BA35BD0",
x"6BA75B77",
x"6BC15B4F",
x"6BE85B59",
x"6C195B92",
x"6C4C5BF6",
x"6C7F5C7A",
x"6CB15D10",
x"6CE55DAE",
x"6D1E5E48",
x"6D655ED2",
x"6DBD5F48",
x"6E285FA5",
x"6EAA5FEA",
x"6F3C601B",
x"6FDE6041",
x"7084605F",
x"712B6080",
x"71C960AB",
x"725B60E0",
x"72D86124",
x"733D6174",
x"738661CB",
x"73AE6224",
x"73B26279",
x"739162C2",
x"734962FD",
x"72DE6324",
x"72536339",
x"71B5633C",
x"7114632F",
x"7081631A",
x"701162FD",
x"6FD462E0",
x"6FD562C4",
x"701E62AB",
x"70AB6298",
x"7172628A",
x"72616283",
x"735F6281",
x"74556286",
x"752D628D",
x"75CF6298",
x"763462A7",
x"765562B4",
x"763562BE",
x"75E262C2",
x"756962BE",
x"74DE62AE",
x"74516290",
x"73D36266",
x"7370622F",
x"732B61F2",
x"730761B2",
x"72FF6176",
x"730A6143",
x"7320611F",
x"7334610D",
x"733B610A",
x"732B6115",
x"72FF6128",
x"72AE613B",
x"723A6145",
x"719E6141",
x"70DE6128",
x"6FFF60F7",
x"6F0360AE",
x"6DF3604F",
x"6CD65FDC",
x"6BB25F5A",
x"6A8D5ECF",
x"696B5E3D",
x"684C5DA8",
x"67315D0E",
x"66165C6E",
x"64F35BC2",
x"63C15B07",
x"62785A36",
x"6111594D",
x"5F895849",
x"5DE1572B",
x"5C1C55F5",
x"5A4554B0",
x"58705363",
x"56B05218",
x"551A50DB",
x"53CA4FBA",
x"52D14EC1",
x"52404DFB",
x"52214D71",
x"52784D27",
x"533A4D22",
x"545C4D60",
x"55C84DDE",
x"57684E96",
x"59204F7F",
x"5ADC508E",
x"5C8751B7",
x"5E1352EE",
x"5F76542B",
x"60AE555D",
x"61BE567F",
x"62A85788",
x"63765870",
x"642D5933",
x"64CE59CD",
x"655E5A3F",
x"65D95A8B",
x"663E5AB5",
x"66875AC3",
x"66B55AC2",
x"66C45AB9",
x"66B85AB5",
x"66965ABD",
x"666B5AD7",
x"663F5B0A",
x"66245B52",
x"66235BAB",
x"66445C0D",
x"668C5C6D",
x"66F85CC1",
x"677F5CFD",
x"68145D18",
x"68A85D12",
x"69285CE7",
x"69855C9E",
x"69B45C3F",
x"69B25BD3",
x"69805B67",
x"69285B07",
x"68BD5ABC",
x"684F5A90",
x"67F95A85",
x"67CB5A9C",
x"67D65AD7",
x"68245B2F",
x"68B15B9F",
x"69765C22",
x"6A625CB3",
x"6B5F5D4B",
x"6C555DE4",
x"6D2E5E7A",
x"6DD85F08",
x"6E475F8E",
x"6E7C6007",
x"6E7F6074",
x"6E5B60D5",
x"6E276129",
x"6DF96174",
x"6DE261B7",
x"6DF061F0",
x"6E2A6222",
x"6E8F624B",
x"6F106266",
x"6FA36274",
x"70346273",
x"70B1625F",
x"710E6239",
x"71476206",
x"715861C8",
x"714C6187",
x"712E6149",
x"710C6117",
x"70F660F3",
x"70F660E0",
x"711160DA",
x"714860DA",
x"719060D9",
x"71DF60C6",
x"72266098",
x"72556046",
x"72625FCC",
x"72425F2B",
x"71F65E6D",
x"71825DA2",
x"70ED5CDF",
x"70485C36",
x"6FA05BC0",
x"6F065B8B",
x"6E845B9F",
x"6E275BFB",
x"6DF05C94",
x"6DE25D59",
x"6DF65E2F",
x"6E245EFE",
x"6E635FAC",
x"6EA46025",
x"6EDF605D",
x"6F076052",
x"6F146008",
x"6F035F91",
x"6ED15EFE",
x"6E7F5E69",
x"6E0F5DE3",
x"6D895D7E",
x"6CF05D42",
x"6C4E5D32",
x"6BA75D46",
x"6AFF5D70",
x"6A545D9F",
x"69A75DBF",
x"68F35DBF",
x"68305D8D",
x"67585D22",
x"66665C7D",
x"65555BA2",
x"64285A9E",
x"62E35982",
x"61945864",
x"604B575A",
x"5F1A5677",
x"5E1655CA",
x"5D515560",
x"5CDC553C",
x"5CC1555E",
x"5D0055BD",
x"5D99564D",
x"5E7D5701",
x"5FA357CA",
x"60F9589A",
x"62705966",
x"63FF5A28",
x"65995ADF",
x"673B5B8D",
x"68E55C35",
x"6A965CE0",
x"6C535D97",
x"6E1E5E5F",
x"6FFD5F3F",
x"71F2603C",
x"73FD6158",
x"76236291",
x"786263E8",
x"7ABB6558",
x"7D2E66DE",
x"7FB8686F",
x"82536A09",
x"84FA6B9E",
x"879E6D27",
x"8A316E9A",
x"8CA16FEE",
x"8EDA7119",
x"90CF7215",
x"926F72DE",
x"93B47376",
x"949873DF",
x"95257420",
x"9563743E",
x"95627446",
x"9532743B",
x"94E7742A",
x"94917416",
x"943C7405",
x"93F373F8",
x"93BB73EF",
x"939873EB",
x"938A73EA",
x"939273EB",
x"93B273EC",
x"93E973EE",
x"943673EE",
x"949C73EE",
x"951873EB",
x"95A573E5",
x"963C73DB",
x"96D773CA",
x"976973B1",
x"97E9738F",
x"984C7365",
x"988A7333",
x"98A172FC",
x"988F72C4",
x"9859728D",
x"98057261",
x"979E7240",
x"972C722F",
x"96BB7231",
x"96537248",
x"95FC7272",
x"95B872AD",
x"958D72F5",
x"957A7344",
x"95807396",
x"959C73EA",
x"95D07437",
x"96177480",
x"966D74C4",
x"96CB74FF",
x"972B7534",
x"97817562",
x"97C37589",
x"97E675A6",
x"97DF75B7",
x"97A875BA",
x"973E75AC",
x"96A5758B",
x"95E47554",
x"950B7509",
x"942C74AC",
x"9356743D",
x"929D73BE",
x"920D7337",
x"91AB72A9",
x"91777217",
x"916C7188",
x"917A7100",
x"91957083",
x"91AE701A",
x"91B66FCB",
x"91A86F9C",
x"91856F93",
x"91586FB5",
x"912E7005",
x"911B707F",
x"9138711F",
x"919571DF",
x"923F72B3",
x"933B738D",
x"94817464",
x"9601752C",
x"979F75DA",
x"993B766C",
x"9AB476DE",
x"9BE97731",
x"9CC2776A",
x"9D31778B",
x"9D35779C",
x"9CD777A3",
x"9C2C77A0",
x"9B4C7798",
x"9A4F7786",
x"994A7767",
x"984A7733",
x"974B76DE",
x"963B765D",
x"9500759D",
x"93747490",
x"9174732D",
x"8EE37168",
x"8BAE6F41",
x"87DC6CC2",
x"83896A00",
x"7EE36719",
x"7A346431",
x"75C96177",
x"71F95F1A",
x"6F095D43",
x"6D345C12",
x"6C945B9B",
x"6D2A5BE0",
x"6ED65CD5",
x"71625E5A",
x"74806049",
x"77E26272",
x"7B3964A1",
x"7E4566AD",
x"80D96876",
x"82DF69E6",
x"845A6AF7",
x"85626BB4",
x"86176C2A",
x"86A76C75",
x"87386CAD",
x"87ED6CEE",
x"88D96D48",
x"8A046DCB",
x"8B6A6E7A",
x"8CFB6F54",
x"8EA4704F",
x"904D715F",
x"91E77279",
x"9360738F",
x"94B27495",
x"95D77582",
x"96D27651",
x"97A176FE",
x"98497786",
x"98CC77EB",
x"9929782C",
x"9963784B",
x"99797850",
x"996D783D",
x"99437818",
x"990377E8",
x"98B477B4",
x"985D777F",
x"9807774B",
x"97B8771B",
x"976E76E8",
x"972976AD",
x"96E07664",
x"968A7603",
x"961E7586",
x"959474E8",
x"94E9742C",
x"941E7357",
x"933B7274",
x"924C7190",
x"916270BE",
x"9091700D",
x"8FE96F8A",
x"8F7C6F40",
x"8F526F30",
x"8F726F58",
x"8FD66FB3",
x"90777034",
x"914870CD",
x"9231716F",
x"9321720D",
x"9400729C",
x"94BB7313",
x"9541736C",
x"958A73A7",
x"959073C4",
x"955A73C7",
x"94F373B3",
x"946C7392",
x"93DD736B",
x"935F7348",
x"930B7334",
x"92F67337",
x"932F7357",
x"93BB7399",
x"949473FE",
x"95AC747E",
x"96EC7512",
x"983375AC",
x"9966763C",
x"9A6076B1",
x"9B0B7702",
x"9B577725",
x"9B3F7713",
x"9AC676D4",
x"9A00766E",
x"990575F1",
x"97F4756C",
x"96E974EF",
x"96017489",
x"954F7444",
x"94E17425",
x"94B9742C",
x"94D07455",
x"951A749A",
x"958474F2",
x"95FA7551",
x"966C75AF",
x"96C87605",
x"9703764A",
x"9717767B",
x"97007692",
x"96C1768C",
x"965A766A",
x"95D37627",
x"952F75C8",
x"94777552",
x"93B174CE",
x"92E47446",
x"921B73C6",
x"9160735A",
x"90B9730D",
x"902E72E8",
x"8FBE72E5",
x"8F6372FE",
x"8F11731F",
x"8EAC732F",
x"8E18730F",
x"8D2E72A1",
x"8BC871C8",
x"89C57072",
x"87116E96",
x"83A76C3D",
x"7F946980",
x"7B026683",
x"76276379",
x"714E6098",
x"6CC95E17",
x"68EC5C21",
x"65FF5AD7",
x"64375A4C",
x"63B45A7A",
x"64765B50",
x"66685CAB",
x"69555E64",
x"6CFC604D",
x"71166241",
x"75566420",
x"798365D5",
x"7D69675E",
x"80F068BB",
x"841169FF",
x"86D56B3A",
x"89526C7C",
x"8B9F6DD4",
x"8DD76F48",
x"900D70D8",
x"9243727B",
x"947B7421",
x"96A775BD",
x"98B4773C",
x"9A8B788D",
x"9C1B79A5",
x"9D5A7A78",
x"9E467B06",
x"9EE97B50",
x"9F537B5A",
x"9FA17B2D",
x"9FF07ADA",
x"A05C7A6E",
x"A0FA79FB",
x"A1DA7996",
x"A2F8794E",
x"A44C7930",
x"A5B57941",
x"A7117981",
x"A83079E3",
x"A8E77A53",
x"A9087ABA",
x"A8757AFC",
x"A71F7AFF",
x"A5087AB3",
x"A2487A11",
x"9F08791D",
x"9B8577F1",
x"97FD76A9",
x"94B1756A",
x"91D9745A",
x"8F9D7395",
x"8E11732F",
x"8D32732A",
x"8CE9737B",
x"8D0A7406",
x"8D6274A9",
x"8DBC7540",
x"8DED75A7",
x"8DD075C7",
x"8D567595",
x"8C817513",
x"8B637450",
x"8A187364",
x"88C5726A",
x"878D717C",
x"868870B1",
x"85CB7016",
x"85566FAB",
x"85246F6C",
x"851E6F4B",
x"852C6F3A",
x"85316F24",
x"85116EFE",
x"84B86EBB",
x"841B6E5B",
x"833B6DDF",
x"82276D4F",
x"80F76CB8",
x"7FD26C2B",
x"7EE36BBA",
x"7E596B76",
x"7E636B6F",
x"7F226BB2",
x"80B46C4B",
x"831F6D3A",
x"865B6E7C",
x"8A467009",
x"8EB771CF",
x"936973BA",
x"981875B1",
x"9C7B7798",
x"A0507953",
x"A3607ACB",
x"A5887BF1",
x"A6BA7CB6",
x"A6FE7D19",
x"A6707D1E",
x"A53B7CCD",
x"A3957C39",
x"A1BB7B75",
x"9FE37A98",
x"9E3D79B7",
x"9CEE78E7",
x"9C0A7837",
x"9B9477B2",
x"9B80775A",
x"9BB6772F",
x"9C157725",
x"9C74772C",
x"9CB17734",
x"9CA87729",
x"9C4576F5",
x"9B7A7689",
x"9A4575E0",
x"98B474F1",
x"96D573C6",
x"94BF7268",
x"928770E5",
x"903C6F4F",
x"8DE36DB3",
x"8B776C1C",
x"88EC6A8D",
x"862C6906",
x"83246781",
x"7FBF65F5",
x"7BFA6456",
x"77D9629F",
x"737860D2",
x"6EFF5EF4",
x"6AA75D14",
x"66AE5B47",
x"635759A9",
x"60D65854",
x"5F59575D",
x"5EF356D9",
x"5FA156CF",
x"614A573D",
x"63C4581B",
x"66D55953",
x"6A3F5ACF",
x"6DCB5C73",
x"71475E24",
x"74905FCC",
x"7798615C",
x"7A6062C8",
x"7CF66410",
x"7F726538",
x"81EC6649",
x"84806753",
x"873F6860",
x"8A2E6980",
x"8D4B6ABB",
x"90846C17",
x"93C26D93",
x"96E46F2D",
x"99CF70D8",
x"9C667288",
x"9E94742C",
x"A04F75B3",
x"A197770D",
x"A274782F",
x"A2FB790F",
x"A34279AC",
x"A3647A08",
x"A37B7A2F",
x"A39C7A2A",
x"A3D77A0E",
x"A43279E7",
x"A4AE79C9",
x"A54279BA",
x"A5E179C4",
x"A67D79E7",
x"A7017A1B",
x"A7617A57",
x"A7917A8E",
x"A78A7AB4",
x"A74A7ABD",
x"A6DA7AA2",
x"A6407A63",
x"A58D7A03",
x"A4CD798E",
x"A4117912",
x"A36778A0",
x"A2D97848",
x"A2707818",
x"A22E7813",
x"A20E783C",
x"A20E788B",
x"A22478F4",
x"A2427965",
x"A26079D0",
x"A2737A23",
x"A2767A54",
x"A2667A61",
x"A2497A4B",
x"A2297A1F",
x"A21179EA",
x"A21179BD",
x"A23979AA",
x"A29779C1",
x"A3327A08",
x"A40E7A7F",
x"A5257B23",
x"A66A7BE5",
x"A7C97CB4",
x"A92B7D7F",
x"AA777E35",
x"AB947EC6",
x"AC6B7F2B",
x"ACF07F61",
x"AD187F6B",
x"ACE77F50",
x"AC637F18",
x"AB9B7ECD",
x"AAA67E78",
x"A99B7E1F",
x"A8927DC6",
x"A7A27D6E",
x"A6DD7D18",
x"A6507CC3",
x"A5FE7C6F",
x"A5E37C1C",
x"A5F67BCC",
x"A6237B7E",
x"A6597B37",
x"A67E7AF9",
x"A6817AC1",
x"A6507A91",
x"A5E47A64",
x"A53B7A39",
x"A45A7A0B",
x"A35379D8",
x"A23979A2",
x"A11F7965",
x"A01C7928",
x"9F3C78EA",
x"9E8A78AF",
x"9E037875",
x"9D9F783E",
x"9D4F7806",
x"9CFE77C6",
x"9C987779",
x"9C08771B",
x"9B3E76A2",
x"9A31760F",
x"98DC755E",
x"9740748D",
x"9566739C",
x"9352728C",
x"910D715A",
x"8EA17006",
x"8C106E8D",
x"89636CF3",
x"86A16B3D",
x"83D36973",
x"810A67A8",
x"7E5D65F5",
x"7BEA6476",
x"79D8634E",
x"78496298",
x"77666270",
x"774F62E2",
x"781863EF",
x"79C96587",
x"7C596791",
x"7FAE69E8",
x"839E6C5E",
x"87F76ECD",
x"8C867110",
x"91147313",
x"957B74D1",
x"99A17651",
x"9D7B77A9",
x"A11778F7",
x"A48D7A60",
x"A8017BFF",
x"AB9F7DED",
x"AF88802F",
x"B3DA82C5",
x"B89B8599",
x"BDBF888E",
x"C3268B7E",
x"C89C8E45",
x"CDE490BC",
x"D2BC92C9",
x"D6E4945B",
x"DA2C9569",
x"DC7595FA",
x"DDB79621",
x"DE0595F5",
x"DD859591",
x"DC6F951B",
x"DB0994B1",
x"D998946F",
x"D85F946C",
x"D79694B8",
x"D7629559",
x"D7D7964C",
x"D8EF9780",
x"DA9998DF",
x"DCAD9A4A",
x"DEFE9B9D",
x"E1549CB6",
x"E37C9D76",
x"E5479DCA",
x"E68F9DA6",
x"E7409D10",
x"E74F9C1F",
x"E6C79AEF",
x"E5BB99AB",
x"E44D987F",
x"E2A19793",
x"E0DF9703",
x"DF2D96E0",
x"DDA9972A",
x"DC6497CE",
x"DB6B98AE",
x"DABB99A3",
x"DA4A9A82",
x"DA059B27",
x"D9D79B76",
x"D9A49B62",
x"D95B9AEC",
x"D8E89A23",
x"D83C991F",
x"D75297FC",
x"D62D96DB",
x"D4D595D2",
x"D35A94F5",
x"D1D3944B",
x"D05793D3",
x"CEFF9384",
x"CDE29355",
x"CD139334",
x"CC999318",
x"CC7492F9",
x"CC9592CE",
x"CCE89297",
x"CD519256",
x"CDAD920A",
x"CDE091B8",
x"CDCE915F",
x"CD6B9100",
x"CCAF909D",
x"CBA59034",
x"CA5A8FC5",
x"C8E78F52",
x"C7628EDC",
x"C5E58E65",
x"C47C8DEF",
x"C3308D7A",
x"C1FF8D04",
x"C0E18C8B",
x"BFCD8C08",
x"BEB68B7A",
x"BD948ADA",
x"BC678A28",
x"BB338964",
x"BA088898",
x"B8FA87CF",
x"B81E8717",
x"B78F8684",
x"B763862B",
x"B7AC861F",
x"B8758671",
x"B9BF872B",
x"BB858853",
x"BDB789E3",
x"C0408BCC",
x"C3028DFA",
x"C5DD904E",
x"C8B092A4",
x"CB5D94D8",
x"CDCA96CA",
x"CFE29858",
x"D198996C",
x"D2DF99F9",
x"D3B499F6",
x"D40B9966",
x"D3D4984F",
x"D2FE96BD",
x"D16A94B5",
x"CEF19244",
x"CB6D8F69",
x"C6B78C28",
x"C0B7887E",
x"B96A8470",
x"B0E48001",
x"A75E7B43",
x"9D29764D",
x"92B87143",
x"888A6C55",
x"7F2267B7",
x"76FC639D",
x"707A6038",
x"6BDE5DAE",
x"693E5C15",
x"688A5B74",
x"698C5BBD",
x"6BED5CD3",
x"6F4F5E8D",
x"734860BF",
x"77796337",
x"7B9665C9",
x"7F6A6858",
x"82DC6AC7",
x"85E36D0C",
x"888E6F20",
x"8AF17108",
x"8D2772C8",
x"8F467465",
x"915D75E1",
x"9373773C",
x"95867872",
x"978E797E",
x"99817A58",
x"9B537AFC",
x"9D007B6A",
x"9E817BA0",
x"9FD97BA8",
x"A10A7B86",
x"A21B7B4A",
x"A3107AF9",
x"A3E97AA2",
x"A4A57A47",
x"A53F79EE",
x"A5B17998",
x"A5F37944",
x"A60078F2",
x"A5D478A3",
x"A5787857",
x"A4F37812",
x"A44D77D8",
x"A39B77B2",
x"A2E677A2",
x"A23B77AA",
x"A19F77CE",
x"A1177809",
x"A09C7856",
x"A02B78AA",
x"9FBC78FC",
x"9F4C7943",
x"9ED47977",
x"9E5A7992",
x"9DE37993",
x"9D76797C",
x"9D1C7951",
x"9CDD7918",
x"9CB978D4",
x"9CA97889",
x"9CA47839",
x"9C9777E1",
x"9C707781",
x"9C1E7716",
x"9B9576A2",
x"9AD27625",
x"99DA75A3",
x"98BF7525",
x"979A74B6",
x"968B7461",
x"95B37430",
x"952E7429",
x"95117450",
x"956674A1",
x"96257516",
x"974075A2",
x"989A7636",
x"9A0D76C1",
x"9B747736",
x"9CAB7788",
x"9D9477B2",
x"9E1877AD",
x"9E2E777E",
x"9DD6772A",
x"9D1C76BA",
x"9C127636",
x"9ACF75AA",
x"99697521",
x"97F974A3",
x"96917436",
x"954173DE",
x"9411739C",
x"93047371",
x"921E7355",
x"915A7344",
x"90B67336",
x"90317321",
x"8FC37302",
x"8F7272CE",
x"8F3B7288",
x"8F227230",
x"8F2B71CB",
x"8F567166",
x"8FA57109",
x"901470C0",
x"909E7090",
x"91397080",
x"91D5708D",
x"926270B1",
x"92CD70E1",
x"93047110",
x"92FA7134",
x"92A77141",
x"92057131",
x"911D7105",
x"8FF970BE",
x"8EAB7066",
x"8D457002",
x"8BD96F97",
x"8A706F29",
x"89106EB1",
x"87AE6E29",
x"863E6D82",
x"84A56CAE",
x"82CB6BA0",
x"80966A51",
x"7DF968BC",
x"7AF366EF",
x"779364F9",
x"73FA62F0",
x"705860F7",
x"6CE95F2B",
x"69EB5DAB",
x"67965C8E",
x"66195BE6",
x"658F5BB8",
x"65FF5C01",
x"67585CB9",
x"69775DCB",
x"6C2D5F24",
x"6F3C60AD",
x"72706250",
x"759763FD",
x"788965A3",
x"7B2F6737",
x"7D8168B1",
x"7F7F6A0F",
x"81356B4B",
x"82B46C66",
x"840D6D62",
x"85526E3F",
x"86906F02",
x"87CF6FAD",
x"891A7044",
x"8A7070CF",
x"8BD87154",
x"8D4C71D7",
x"8ED0725C",
x"905F72E8",
x"91F1737B",
x"937E7416",
x"94FA74B9",
x"9656755B",
x"978375FC",
x"98747696",
x"991F7720",
x"99807795",
x"999777F1",
x"996F782A",
x"9911783E",
x"98917829",
x"980077E8",
x"976E777C",
x"96E976E7",
x"96787630",
x"96257564",
x"95ED7490",
x"95D273C4",
x"95D37313",
x"95F07290",
x"962B7248",
x"96877247",
x"970D7290",
x"97BF7325",
x"98A173F9",
x"99B57501",
x"9AF37627",
x"9C52775A",
x"9DC27881",
x"9F2C798B",
x"A07D7A68",
x"A19F7B11",
x"A27E7B7E",
x"A30C7BB3",
x"A3427BB3",
x"A31B7B86",
x"A29E7B36",
x"A1D37ACA",
x"A0C37A4B",
x"9F8079C0",
x"9E17792C",
x"9C947896",
x"9B087803",
x"997E7779",
x"980376FE",
x"96A27697",
x"9566764E",
x"94597625",
x"9383761C",
x"92EA7631",
x"92907661",
x"9274769B",
x"929376D4",
x"92DF76FC",
x"934D7705",
x"93CF76E5",
x"94537696",
x"94C9761A",
x"95227578",
x"955274BB",
x"954C73F5",
x"950A7336",
x"9488728F",
x"93CC720A",
x"92D971B0",
x"91BF7183",
x"908B717E",
x"8F587199",
x"8E3971CA",
x"8D4D720A",
x"8CA87251",
x"8C5C7299",
x"8C7472DF",
x"8CF07326",
x"8DC57371",
x"8ED973BE",
x"90107410",
x"91467465",
x"925974B7",
x"932A7501",
x"93A27534",
x"93B8754B",
x"936F753D",
x"92D57505",
x"91FD74A0",
x"91037416",
x"8FFC736C",
x"8EF972AF",
x"8E0471E9",
x"8D1B7127",
x"8C31706C",
x"8B356FBB",
x"8A116F0F",
x"88AE6E5B",
x"86FE6D92",
x"84FB6CA1",
x"82A56B7C",
x"800C6A19",
x"7D446876",
x"7A6C66A1",
x"77A864AF",
x"751D62BE",
x"72E960F4",
x"712E5F78",
x"70035E70",
x"6F795DF6",
x"6F9A5E18",
x"70665ED6",
x"71D86022",
x"73E261DF",
x"766F63E6",
x"79666613",
x"7CAE683C",
x"80286A48",
x"83B86C26",
x"87456DD1",
x"8ABE6F52",
x"8E1070BE",
x"9138722A",
x"943273AD",
x"97047558",
x"99B47733",
x"9C49793D",
x"9ECD7B67",
x"A14A7D9C",
x"A3C27FC2",
x"A63681C2",
x"A8A28381",
x"AB0084F4",
x"AD428612",
x"AF5A86DD",
x"B136875C",
x"B2C28799",
x"B3ED87A7",
x"B4A5878D",
x"B4DE8756",
x"B4978704",
x"B3D0869B",
x"B2978617",
x"B0FE8576",
x"AF2284B5",
x"AD1F83D4",
x"AB1882DC",
x"A92581D0",
x"A75E80BD",
x"A5D47FB0",
x"A48D7EB9",
x"A38A7DE3",
x"A2C37D37",
x"A2357CC1",
x"A1D67C84",
x"A1A27C7F",
x"A19A7CAF",
x"A1BF7D0E",
x"A2187D94",
x"A2A97E32",
x"A3767EDD",
x"A4737F84",
x"A594801B",
x"A6C08091",
x"A7D980D9",
x"A8BA80E8",
x"A94580B7",
x"A9608049",
x"A9007F9F",
x"A8297ECA",
x"A6F07DDD",
x"A57D7CF1",
x"A4027C22",
x"A2BB7B8E",
x"A1DD7B4D",
x"A19B7B71",
x"A2117C05",
x"A34C7D02",
x"A53D7E5D",
x"A7C27FF7",
x"AAA281B0",
x"AD9B8363",
x"B06A84E6",
x"B2C78615",
x"B47F86DC",
x"B56D8729",
x"B5828700",
x"B4C78669",
x"B35C857D",
x"B16B845A",
x"AF2C8321",
x"ACD981F1",
x"AAA380E6",
x"A8B9800F",
x"A7367F7A",
x"A6297F23",
x"A5917F08",
x"A5647F19",
x"A58F7F4A",
x"A5FA7F8E",
x"A68D7FD9",
x"A7368020",
x"A7E98064",
x"A89A809F",
x"A94580D6",
x"A9E98107",
x"AA878136",
x"AB1C8163",
x"ABA8818C",
x"AC2381AD",
x"AC8881C3",
x"ACCC81C7",
x"ACE681B0",
x"ACCF817A",
x"AC80811F",
x"ABF7809C",
x"AB367FF0",
x"AA467F1E",
x"A92B7E2D",
x"A7F37D22",
x"A6A67C05",
x"A54C7AE4",
x"A3E679C4",
x"A27078AA",
x"A0DF7799",
x"9F1D768B",
x"9D107572",
x"9A9A7444",
x"979E72EB",
x"94037155",
x"8FBC6F75",
x"8ACF6D44",
x"85506AC4",
x"7F6D6800",
x"79626513",
x"737C621A",
x"6E0F5F41",
x"696D5CAE",
x"65DF5A87",
x"639758EE",
x"62B057F5",
x"632657A4",
x"64D757F5",
x"678A58D6",
x"6AF55A2E",
x"6EC55BDA",
x"72AB5DBB",
x"76655FB1",
x"79C261A2",
x"7CAB637D",
x"7F1B6538",
x"812566D2",
x"82E6684C",
x"848169AE",
x"861B6B03",
x"87CD6C51",
x"89AB6D9D",
x"8BB86EEE",
x"8DF17043",
x"904B719C",
x"92B672F6",
x"9527744E",
x"979175A3",
x"99F076F2",
x"9C42783C",
x"9E88797E",
x"A0C67AB9",
x"A2F87BEB",
x"A5197D14",
x"A7217E2F",
x"A9007F37",
x"AAA5802B",
x"ABFE8100",
x"ACFF81B0",
x"ADA28237",
x"ADE78292",
x"ADD482BD",
x"AD7B82BC",
x"ACF1828F",
x"AC49823D",
x"AB9781CF",
x"AAED814C",
x"AA5680BD",
x"A9D9802D",
x"A9737FA2",
x"A9217F23",
x"A8D97EB7",
x"A8957E61",
x"A84F7E20",
x"A8017DF7",
x"A7AB7DE1",
x"A74F7DDD",
x"A6EE7DE5",
x"A68E7DF1",
x"A62E7DF8",
x"A5CD7DF1",
x"A56A7DD3",
x"A4FD7D96",
x"A4807D37",
x"A3EE7CB4",
x"A3467C13",
x"A28B7B5B",
x"A1C87A9D",
x"A10D79EE",
x"A0707961",
x"A008790F",
x"9FEC7908",
x"A02C795A",
x"A0CD7A09",
x"A1CA7B0F",
x"A3127C5A",
x"A4847DD1",
x"A5FD7F54",
x"A75080C2",
x"A85D81F8",
x"A90482DE",
x"A9388360",
x"A8F8837B",
x"A8568335",
x"A76D829F",
x"A66481D3",
x"A56280EB",
x"A4878005",
x"A3EC7F36",
x"A39A7E8E",
x"A38B7E11",
x"A3AE7DB9",
x"A3E67D7E",
x"A4177D50",
x"A4217D1F",
x"A3F47CDE",
x"A3847C86",
x"A2D77C18",
x"A1FE7B99",
x"A1147B18",
x"A03B7AA2",
x"9F917A4B",
x"9F357A23",
x"9F407A33",
x"9FBE7A81",
x"A0B07B0C",
x"A2127BCE",
x"A3D67CBC",
x"A5E77DC6",
x"A82F7EDD",
x"AA977FF0",
x"AD0780F5",
x"AF6981E0",
x"B1AC82A9",
x"B3BD834F",
x"B58C83CC",
x"B70C8423",
x"B82C8452",
x"B8DB8459",
x"B90B8433",
x"B8A683DC",
x"B7998347",
x"B5CD826D",
x"B32F813F",
x"AFAE7FAF",
x"AB437DB7",
x"A5EB7B4E",
x"9FB97879",
x"98CC7543",
x"915671C0",
x"899A6E0F",
x"81E56A52",
x"7A9166B8",
x"73F86369",
x"6E686090",
x"6A265E4F",
x"675F5CBC",
x"662A5BE9",
x"667D5BD0",
x"68385C6A",
x"6B265D9E",
x"6EFF5F4D",
x"73756155",
x"783C6390",
x"7D1165DB",
x"81BB6819",
x"86146A34",
x"8A0A6C20",
x"8D9B6DD8",
x"90D06F5F",
x"93BB70BE",
x"96717203",
x"9904733A",
x"9B80746F",
x"9DE475A9",
x"A02976E8",
x"A2427827",
x"A418795E",
x"A59B7A81",
x"A6BA7B82",
x"A7757C5A",
x"A7D27D08",
x"A7E37D8E",
x"A7C67DF8",
x"A7A27E59",
x"A7977EC4",
x"A7C27F4D",
x"A8388002",
x"A8F880EA",
x"A9F681FB",
x"AB158329",
x"AC2F8457",
x"AD178568",
x"ADAC863C",
x"ADD286B8",
x"AD7D86C9",
x"ACB6866C",
x"AB9285A7",
x"AA39848F",
x"A8D38342",
x"A78D81E0",
x"A688808C",
x"A5DC7F63",
x"A58E7E77",
x"A5977DD1",
x"A5E07D6F",
x"A64F7D49",
x"A6C37D4A",
x"A7247D61",
x"A7597D7B",
x"A75A7D87",
x"A7267D7B",
x"A6C57D54",
x"A6427D15",
x"A5AE7CC3",
x"A5157C6A",
x"A4817C13",
x"A3F77BCA",
x"A37A7B96",
x"A3057B7E",
x"A2977B81",
x"A2287B9F",
x"A1B37BD3",
x"A13B7C16",
x"A0BC7C63",
x"A03B7CAD",
x"9FBE7CEE",
x"9F487D1F",
x"9EDD7D39",
x"9E817D36",
x"9E367D15",
x"9DF87CD3",
x"9DC67C72",
x"9D987BF5",
x"9D697B64",
x"9D2F7AC4",
x"9CE47A1F",
x"9C86797F",
x"9C1078EE",
x"9B837874",
x"9AE37816",
x"9A3977D4",
x"998B77AA",
x"98E27793",
x"98437782",
x"97B57768",
x"97367737",
x"96C576E7",
x"965F766F",
x"95FE75D0",
x"95A57512",
x"95527444",
x"950B7378",
x"94DA72C5",
x"94CC7243",
x"94EC7200",
x"95427208",
x"95D5725B",
x"969E72F4",
x"979473BE",
x"98A274A7",
x"99B17597",
x"9AA87675",
x"9B73772F",
x"9C0177B7",
x"9C4F780C",
x"9C61782F",
x"9C487829",
x"9C147805",
x"9BD677D0",
x"9B9C7792",
x"9B67774A",
x"9B2876F5",
x"9AC67686",
x"9A1B75F1",
x"98FA7520",
x"973B7408",
x"94C1729F",
x"917E70E4",
x"8D836EE2",
x"88F36CAD",
x"840D6A65",
x"7F24682D",
x"7A90662B",
x"76AB6483",
x"73C26352",
x"720C62AE",
x"719E629D",
x"7279631B",
x"7474641B",
x"77586586",
x"7AD8673E",
x"7EA46924",
x"82746B1D",
x"86096D0F",
x"89376EE5",
x"8BE67094",
x"8E187217",
x"8FD8736B",
x"913E7495",
x"92697595",
x"93737674",
x"94717733",
x"957477D7",
x"96817861",
x"979778D0",
x"98B27926",
x"99C87961",
x"9AD37985",
x"9BCC7990",
x"9CAF7986",
x"9D7A796B",
x"9E2B793E",
x"9EC07906",
x"9F3978C3",
x"9F917879",
x"9FC2782A",
x"9FCC77D8",
x"9FAB7786",
x"9F62773A",
x"9EF776F4",
x"9E7476BA",
x"9DE6768F",
x"9D597678",
x"9CDD7675",
x"9C7A7686",
x"9C3676AD",
x"9C1576E2",
x"9C107726",
x"9C1F776F",
x"9C3977BC",
x"9C4F7805",
x"9C567848",
x"9C467882",
x"9C1578B0",
x"9BC278D0",
x"9B4878DE",
x"9AA878DA",
x"99E478BA",
x"98FB787E",
x"97F0781C",
x"96C37792",
x"957B76DE",
x"941B7602",
x"92AC7503",
x"913B73EE",
x"8FCF72D0",
x"8E7A71BA",
x"8D4870C0",
x"8C436FF2",
x"8B746F5B",
x"8AE26F00",
x"8A876EE1",
x"8A5F6EF6",
x"8A636F2E",
x"8A846F7A",
x"8AB86FC4",
x"8AEF6FFA",
x"8B1F700F",
x"8B426FF9",
x"8B506FB7",
x"8B496F4E",
x"8B2E6ECA",
x"8B046E3A",
x"8AD26DB0",
x"8A9E6D3B",
x"8A6F6CEB",
x"8A4B6CC7",
x"8A346CD2",
x"8A296D0C",
x"8A2B6D68",
x"8A316DD9",
x"8A356E52",
x"8A2F6EC3",
x"8A1A6F1A",
x"89F26F4F",
x"89B46F5E",
x"89666F47",
x"89146F12",
x"88C66ECB",
x"88906E80",
x"887C6E44",
x"88976E24",
x"88EA6E2A",
x"89736E5B",
x"8A2C6EB5",
x"8B066F30",
x"8BEA6FBD",
x"8CBF704A",
x"8D6A70C3",
x"8DD27117",
x"8DE5713B",
x"8D977126",
x"8CE970D7",
x"8BE57054",
x"8A9D6FA6",
x"892D6EDC",
x"87AE6E03",
x"863E6D24",
x"84F06C48",
x"83CF6B6F",
x"82D86A96",
x"81FC69B1",
x"812168B4",
x"80226790",
x"7EDC6638",
x"7D2B64A7",
x"7AFE62DA",
x"784E60DD",
x"752D5EBD",
x"71BE5C97",
x"6E3B5A8A",
x"6AE858B6",
x"68105742",
x"65F85649",
x"64D455E0",
x"64C95615",
x"65DE56E4",
x"67FF5843",
x"6B025A1B",
x"6EA75C4C",
x"72AA5EB3",
x"76C2612E",
x"7AB26398",
x"7E4965DB",
x"816D67DF",
x"8414699A",
x"86496B09",
x"88256C33",
x"89C66D1E",
x"8B4E6DDF",
x"8CDA6E86",
x"8E816F29",
x"90506FD8",
x"924A70AA",
x"946D71A9",
x"96AE72DF",
x"98FB744D",
x"9B4875EC",
x"9D7E77AF",
x"9F8F797C",
x"A16B7B39",
x"A3027CC7",
x"A44D7E07",
x"A5407EE0",
x"A5DA7F3D",
x"A6197F20",
x"A6077E91",
x"A5AB7DA2",
x"A5157C78",
x"A4567B3A",
x"A3807A11",
x"A2A27922",
x"A1D0788B",
x"A114785B",
x"A07A7893",
x"A0077929",
x"9FC27A02",
x"9FAB7B01",
x"9FC37C02",
x"A00A7CE5",
x"A07B7D92",
x"A1127DF5",
x"A1C57E08",
x"A2877DD0",
x"A3497D56",
x"A3FB7CAD",
x"A48B7BEA",
x"A4EC7B1F",
x"A50F7A61",
x"A4F479BD",
x"A49C7940",
x"A41178EB",
x"A36078C0",
x"A29B78B6",
x"A1D778C6",
x"A12478E2",
x"A09278FE",
x"A02B7910",
x"9FF4790E",
x"9FF378F5",
x"A02278C4",
x"A0807883",
x"A107783D",
x"A1B277FC",
x"A27777D1",
x"A34F77C7",
x"A42F77E8",
x"A50D7836",
x"A5D778AF",
x"A6877947",
x"A70B79F4",
x"A75C7AA2",
x"A7717B3E",
x"A74C7BBD",
x"A6ED7C0E",
x"A6597C29",
x"A59B7C0C",
x"A4BB7BBA",
x"A3BD7B36",
x"A2AB7A86",
x"A18579B3",
x"A04C78C6",
x"9EFE77C6",
x"9D9F76BC",
x"9C2F75AF",
x"9AB674A9",
x"994273B3",
x"97DF72DB",
x"96A2722B",
x"959F71AD",
x"94E4716B",
x"947E7166",
x"947171A4",
x"94B9721C",
x"954C72C4",
x"96147390",
x"96FB746F",
x"97E6754D",
x"98BC7619",
x"996476C4",
x"99CF7743",
x"99F3778F",
x"99CF77A5",
x"99697786",
x"98CD773A",
x"981176CA",
x"9748763C",
x"96807599",
x"95C874E8",
x"95217429",
x"9487735E",
x"93E67280",
x"93247188",
x"921E706E",
x"90B26F27",
x"8EC16DAE",
x"8C366C03",
x"890D6A26",
x"85536821",
x"812E6606",
x"7CCE63E9",
x"787661E4",
x"74706015",
x"71015E95",
x"6E685D7D",
x"6CCE5CDF",
x"6C495CC3",
x"6CD95D2E",
x"6E635E18",
x"70BB5F74",
x"73A7612F",
x"76EC632F",
x"7A4C655C",
x"7D9A679B",
x"80B169D8",
x"837F6BFD",
x"86016DFD",
x"88466FCF",
x"8A62716F",
x"8C7172DC",
x"8E90741A",
x"90D37530",
x"934F7625",
x"960A76FF",
x"98FD77C8",
x"9C1E7889",
x"9F547947",
x"A2857A09",
x"A5927AD4",
x"A85D7BAA",
x"AAC97C91",
x"ACC37D84",
x"AE3D7E81",
x"AF387F82",
x"AFB9807C",
x"AFCD8164",
x"AF8C8229",
x"AF0C82BC",
x"AE64830C",
x"ADAB8311",
x"ACF182C3",
x"AC3B8223",
x"AB8F813B",
x"AAEB8019",
x"AA4D7ED7",
x"A9AF7D8E",
x"A9157C5B",
x"A8817B5D",
x"A7FD7AA9",
x"A7987A51",
x"A75E7A5B",
x"A7617AC4",
x"A7A87B84",
x"A8357C82",
x"A9057DA8",
x"AA087ED7",
x"AB287FF2",
x"AC4780E6",
x"AD488196",
x"AE0F81F7",
x"AE888202",
x"AEA481B7",
x"AE5E8121",
x"ADC2804C",
x"ACE37F4C",
x"ABDD7E3D",
x"AAD07D35",
x"A9E37C4A",
x"A9327B95",
x"A8DA7B25",
x"A8EA7B01",
x"A9667B2D",
x"AA497BA3",
x"AB827C5B",
x"ACFB7D41",
x"AE997E47",
x"B0467F59",
x"B1E78068",
x"B370816A",
x"B4D48254",
x"B6158328",
x"B73283E0",
x"B8338481",
x"B91C850D",
x"B9EE8584",
x"BAA685E6",
x"BB3D8631",
x"BBA8865E",
x"BBDA866D",
x"BBCA8659",
x"BB718622",
x"BAD085CD",
x"B9ED8560",
x"B8D784E1",
x"B7A0845D",
x"B65E83DC",
x"B5258364",
x"B4078300",
x"B30F82AD",
x"B243826E",
x"B1A8823F",
x"B139821F",
x"B0F7820C",
x"B0DB8205",
x"B0E6820B",
x"B10F821C",
x"B154823C",
x"B1B08266",
x"B2188297",
x"B28182C7",
x"B2DD82F1",
x"B322830B",
x"B344830B",
x"B33F82ED",
x"B31282B1",
x"B2C58257",
x"B26181E7",
x"B1F68168",
x"B18780E4",
x"B119805D",
x"B0A27FCF",
x"B00B7F32",
x"AF337E75",
x"ADF17D81",
x"AC217C3F",
x"A99A7A9C",
x"A64C7890",
x"A238761D",
x"9D747354",
x"98317057",
x"92AE6D4E",
x"8D396A70",
x"882567ED",
x"83BB65F3",
x"803964A1",
x"7DC86407",
x"7C796421",
x"7C4664D9",
x"7D1A6610",
x"7EC8679A",
x"8122694C",
x"83F66B03",
x"87106CA4",
x"8A4B6E20",
x"8D866F7C",
x"90AB70C1",
x"93B17206",
x"96947361",
x"995774E5",
x"9C0476A0",
x"9EA47892",
x"A1407AB4",
x"A3E17CF2",
x"A68D7F35",
x"A9458160",
x"AC078359",
x"AEC7850D",
x"B1818670",
x"B422877E",
x"B69C8842",
x"B8DD88C8",
x"BADC8924",
x"BC8E896A",
x"BDEF89AF",
x"BF048A01",
x"BFD38A6A",
x"C0678AEC",
x"C0D08B81",
x"C11C8C22",
x"C1588CC5",
x"C18E8D5C",
x"C1C68DDB",
x"C2018E39",
x"C23F8E70",
x"C27E8E7C",
x"C2B78E5D",
x"C2E88E17",
x"C3098DAC",
x"C3198D25",
x"C3158C87",
x"C2FF8BDC",
x"C2DB8B28",
x"C2B38A79",
x"C28F89D6",
x"C27F894C",
x"C29288E6",
x"C2D888AF",
x"C36388B1",
x"C43788F3",
x"C55D8979",
x"C6CD8A42",
x"C87F8B46",
x"CA608C7E",
x"CC558DDB",
x"CE498F4B",
x"D02290BE",
x"D1D09227",
x"D350937A",
x"D4A294B1",
x"D5D495C8",
x"D6FC96C4",
x"D83097A5",
x"D97F9875",
x"DAF59935",
x"DC8C99E5",
x"DE349A80",
x"DFCE9B02",
x"E1349B5B",
x"E2419B85",
x"E2D09B75",
x"E2CB9B29",
x"E22F9AA3",
x"E10C99F0",
x"DF839920",
x"DDC4984B",
x"DC039786",
x"DA7496E8",
x"D939967C",
x"D8679648",
x"D7F99641",
x"D7D79655",
x"D7D29666",
x"D7B29655",
x"D73995FD",
x"D6369547",
x"D486941E",
x"D21A927D",
x"CEFF9070",
x"CB578E0E",
x"C7578B79",
x"C33D88D9",
x"BF4D8656",
x"BBBD8418",
x"B8B78239",
x"B65080C9",
x"B4857FCC",
x"B33A7F35",
x"B2477EF0",
x"B1727EDB",
x"B0857ED7",
x"AF4D7EC1",
x"ADA57E7B",
x"AB807DF1",
x"A8DD7D19",
x"A5DD7BF4",
x"A2AB7A91",
x"9F7D7903",
x"9C8B7768",
x"9A0775DE",
x"980B747C",
x"96A17354",
x"95B2726C",
x"951471BE",
x"94817133",
x"93AE70AD",
x"924A7005",
x"90146F17",
x"8CE06DC2",
x"889F6BF2",
x"836A69A6",
x"7D7766EB",
x"771B63E2",
x"70BE60BF",
x"6ACF5DB9",
x"65B45B0D",
x"61C058EB",
x"5F26577E",
x"5DFA56D6",
x"5E2D56F5",
x"5F8D57C3",
x"61D4591B",
x"64AE5ACA",
x"67CB5C9C",
x"6ADE5E5F",
x"6DAE5FE7",
x"701A611A",
x"721361E8",
x"739E6255",
x"74D1626C",
x"75C66242",
x"769961F3",
x"775C6195",
x"78206141",
x"78E66103",
x"79A860E7",
x"7A5C60F2",
x"7AF46121",
x"7B666173",
x"7BAB61E4",
x"7BC56273",
x"7BBB631B",
x"7B9D63DD",
x"7B7964BA",
x"7B6065AD",
x"7B6366B7",
x"7B8C67D1",
x"7BDB68F2",
x"7C4F6A0F",
x"7CE66B1A",
x"7D936C06",
x"7E4B6CC2",
x"7F046D45",
x"7FB86D88",
x"80606D83",
x"80FC6D3B",
x"818A6CB7",
x"820D6C03",
x"82866B2D",
x"82F96A45",
x"8363695B",
x"83C4687F",
x"841467BA",
x"844B6713",
x"8463668E",
x"8450662B",
x"841065E5",
x"839E65B7",
x"82FD659A",
x"82326587",
x"814E657A",
x"805D656D",
x"7F76655F",
x"7EA8654F",
x"7E06653F",
x"7D956531",
x"7D596528",
x"7D4E6528",
x"7D636532",
x"7D896548",
x"7DA86566",
x"7DB1658D",
x"7D9565B5",
x"7D5365DE",
x"7CED6600",
x"7C74661A",
x"7BFC6628",
x"7B9E6631",
x"7B736634",
x"7B8C663C",
x"7BF3664F",
x"7CA76675",
x"7D9A66B4",
x"7EB7670E",
x"7FE26783",
x"8100680C",
x"81F9689E",
x"82B96930",
x"833C69B2",
x"83836A1E",
x"83976A6C",
x"838D6A9A",
x"83736AAA",
x"835C6AA1",
x"83526A87",
x"83586A62",
x"836A6A35",
x"837F6A03",
x"838769C9",
x"83736982",
x"83396924",
x"82CF68AD",
x"82356819",
x"816F676B",
x"808666A8",
x"7F8465DE",
x"7E776515",
x"7D69645F",
x"7C5F63C1",
x"7B5C6342",
x"7A6262E0",
x"796A6293",
x"78776250",
x"7784620D",
x"769761BE",
x"75B7615D",
x"74EC60EE",
x"74426076",
x"73C75FFE",
x"73825F97",
x"73725F4B",
x"73945F1E",
x"73D85F0E",
x"74275F11",
x"74605F11",
x"74635EF6",
x"740E5EA2",
x"73445E00",
x"71ED5CFE",
x"70035B9B",
x"6D8759DD",
x"6A9057DD",
x"673B55BD",
x"63B553A5",
x"603051C0",
x"5CE35032",
x"5A004F18",
x"57B64E85",
x"56244E7B",
x"55654EF2",
x"557B4FD7",
x"565F510E",
x"57FE527A",
x"5A3153FE",
x"5CD55584",
x"5FBB56F5",
x"62B45847",
x"65995971",
x"68425A73",
x"6A975B4D",
x"6C865C04",
x"6E045C9A",
x"6F175D12",
x"6FC65D74",
x"70265DC3",
x"70455E06",
x"703C5E3D",
x"701D5E74",
x"6FFA5EAE",
x"6FDF5EF1",
x"6FD15F42",
x"6FD45F9F",
x"6FE5600A",
x"6FFF607C",
x"701E60EE",
x"703F615C",
x"706261BB",
x"70846206",
x"70AE6239",
x"70E36256",
x"712B6260",
x"7189625D",
x"71FF6256",
x"72876252",
x"731A6259",
x"73AD626F",
x"742E6294",
x"749162C6",
x"74CE6300",
x"74DE6339",
x"74C4636D",
x"74896394",
x"743E63AA",
x"73F663AE",
x"73C563A3",
x"73BD638B",
x"73E66372",
x"74456359",
x"74D16348",
x"75796344",
x"7624634E",
x"76BA6363",
x"771D6383",
x"773863A5",
x"76FD63C6",
x"766863E0",
x"757F63EF",
x"745363ED",
x"72FD63DD",
x"719D63BE",
x"704E6391",
x"6F30635A",
x"6E56631D",
x"6DD462DA",
x"6DAB6295",
x"6DDB624F",
x"6E566207",
x"6F0C61BF",
x"6FE36179",
x"70C86135",
x"71A660F4",
x"726860BC",
x"7304608E",
x"7373606D",
x"73B46059",
x"73CB6056",
x"73BE6063",
x"7397607D",
x"735C60A1",
x"731660CC",
x"72C960FC",
x"7279612B",
x"72276159",
x"71D36186",
x"718261AF",
x"713061D9",
x"70E26203",
x"709E622D",
x"70686253",
x"70426273",
x"70326289",
x"7037628B",
x"704C6279",
x"706F624B",
x"70966201",
x"70B761A2",
x"70C96132",
x"70C760BE",
x"70A86055",
x"706F6004",
x"701E5FD9",
x"6FBA5FDA",
x"6F48600A",
x"6ED46063",
x"6E6060D8",
x"6DF36155",
x"6D8C61C3",
x"6D28620E",
x"6CC46224",
x"6C5861F4",
x"6BDE617E",
x"6B4E60C3",
x"6AA65FD5",
x"69DF5EC2",
x"68FD5DA4",
x"68025C90",
x"66F25B97",
x"65D25AC3",
x"64AB5A1B",
x"63875997",
x"626C592C",
x"616558CA",
x"60765861",
x"5FA957E4",
x"5F03574D",
x"5E88569B",
x"5E3855D7",
x"5E1A5515",
x"5E2D546A",
x"5E7253F1",
x"5EE853C4",
x"5F9353F5",
x"60735491",
x"618D5599",
x"62E35707",
x"647558C6",
x"66425ABC",
x"68475CC9",
x"6A795ECD",
x"6CCB60AB",
x"6F2B6249",
x"71846397",
x"73BF648E",
x"75C86531",
x"778A6586",
x"78FD659E",
x"7A1B658E",
x"7AEA6569",
x"7B796542",
x"7BD66527",
x"7C206525",
x"7C696542",
x"7CCB6581",
x"7D5265E0",
x"7E07665C",
x"7EE666ED",
x"7FE3678E",
x"80F0683B",
x"81F468EC",
x"82DF699E",
x"839B6A4B",
x"84216AF0",
x"846F6B8A",
x"848D6C16",
x"84896C90",
x"84776CF5",
x"846C6D41",
x"847A6D76",
x"84B16D92",
x"85146D96",
x"85A46D88",
x"86586D6B",
x"87256D4A",
x"87FD6D2E",
x"88D36D24",
x"89A26D38",
x"8A666D73",
x"8B246DDE",
x"8BE56E7C",
x"8CB46F4A",
x"8D9C7043",
x"8EA77157",
x"8FD37276",
x"911D738C",
x"92797482",
x"93D57547",
x"951C75D0",
x"963B7615",
x"9721761A",
x"97C575EB",
x"98287599",
x"9853753B",
x"985874EB",
x"984F74BD",
x"985474C4",
x"98847509",
x"98F0758F",
x"99A8764E",
x"9AAE7737",
x"9BFB7837",
x"9D7B7937",
x"9F157A25",
x"A0A97AEA",
x"A21A7B7C",
x"A3477BD4",
x"A41F7BF2",
x"A4947BD9",
x"A4A47B92",
x"A4567B28",
x"A3BC7AA8",
x"A2EB7A1C",
x"A1FD7990",
x"A1087909",
x"A024788C",
x"9F5C7818",
x"9EBB77A9",
x"9E3D773C",
x"9DE076C8",
x"9D9A7647",
x"9D5F75B3",
x"9D21750B",
x"9CDA744D",
x"9C847382",
x"9C1C72B4",
x"9BA871F4",
x"9B2E714F",
x"9AB670DB",
x"9A4A70A3",
x"99F070B3",
x"99AC7109",
x"997D71A0",
x"995C7266",
x"99407347",
x"991D7423",
x"98E774DE",
x"9894755C",
x"981E758C",
x"97847561",
x"96CB74D8",
x"95FA73FB",
x"951B72D8",
x"94367185",
x"934B7013",
x"92566E94",
x"91496D14",
x"900D6B96",
x"8E866A16",
x"8C97688D",
x"8A2B66F2",
x"8737653B",
x"83BB6366",
x"7FD3617A",
x"7BA75F84",
x"77725D9B",
x"737C5BDA",
x"700A5A64",
x"6D635953",
x"6BB858C3",
x"6B2A58BF",
x"6BBA594D",
x"6D555A63",
x"6FCE5BF0",
x"72EB5DD6",
x"76655FF4",
x"79F96229",
x"7D6D6458",
x"80966662",
x"83586835",
x"85AF69CC",
x"87AB6B21",
x"89666C3E",
x"8B006D30",
x"8CA16E06",
x"8E696ED7",
x"90706FB0",
x"92C370A6",
x"956371C0",
x"98427305",
x"9B497474",
x"9E5D7603",
x"A15A77A7",
x"A4227950",
x"A6977AEA",
x"A8A47C64",
x"AA387DAF",
x"AB537EC1",
x"ABFA7F94",
x"AC368029",
x"AC1E8084",
x"ABC580AF",
x"AB3D80AF",
x"AA9F8091",
x"A9F48059",
x"A9458008",
x"A8957FA2",
x"A7E17F22",
x"A7227E88",
x"A6547DCF",
x"A5707CF8",
x"A4767C0B",
x"A3677B12",
x"A24F7A1C",
x"A1397937",
x"A0357877",
x"9F5277E7",
x"9E9D7790",
x"9E1C7775",
x"9DD37790",
x"9DBC77D5",
x"9DCC7834",
x"9DF4789B",
x"9E2978F5",
x"9E5F793A",
x"9E887960",
x"9EA77965",
x"9EB97951",
x"9EC6792F",
x"9ED47909",
x"9EE978EB",
x"9F0778DD",
x"9F2878DE",
x"9F4678EB",
x"9F5478FB",
x"9F4378FE",
x"9F0778E8",
x"9E9578B3",
x"9DF07858",
x"9D1F77E0",
x"9C357754",
x"9B4576C8",
x"9A6D7654",
x"99C27608",
x"995A75F4",
x"99407620",
x"99767688",
x"99F1771F",
x"9AA677D2",
x"9B81788B",
x"9C6C792D",
x"9D5579A5",
x"9E2C79E7",
x"9EE979EA",
x"9F8579B4",
x"A0017950",
x"A05C78CA",
x"A0977837",
x"A0AF77A5",
x"A0A4771F",
x"A07376AC",
x"A0177650",
x"9F947609",
x"9EEC75D2",
x"9E2775AC",
x"9D557592",
x"9C847586",
x"9BC8758B",
x"9B3275A2",
x"9AD075D1",
x"9AAE7619",
x"9ACA7678",
x"9B2576EA",
x"9BB17765",
x"9C6177E1",
x"9D25784E",
x"9DEE78A2",
x"9EAE78D6",
x"9F5C78E1",
x"9FF478C8",
x"A077788F",
x"A0EA7841",
x"A15077EA",
x"A1AE7795",
x"A2037750",
x"A246771D",
x"A26676FF",
x"A24C76EB",
x"A1D276D0",
x"A0D3769B",
x"9F28762F",
x"9CAE7574",
x"994F7452",
x"950372BD",
x"8FD870AE",
x"89F36E30",
x"838E6B55",
x"7CF3683F",
x"76766518",
x"706F6210",
x"6B2E5F52",
x"66F65D0B",
x"63F35B59",
x"623A5A4F",
x"61C159F0",
x"62695A35",
x"64035B08",
x"664C5C49",
x"69065DD6",
x"6BEC5F8B",
x"6EC86146",
x"717262EF",
x"73D16470",
x"75DC65C5",
x"779B66EC",
x"791E67E9",
x"7A7E68C8",
x"7BD36997",
x"7D386A62",
x"7EBA6B30",
x"80606C06",
x"822A6CE5",
x"840B6DC7",
x"85F16EA0",
x"87C16F65",
x"89637008",
x"8AC1707C",
x"8BC670BA",
x"8C7070BD",
x"8CBE7088",
x"8CBB7024",
x"8C7E6F9D",
x"8C1E6F06",
x"8BB96E6E",
x"8B676DE3",
x"8B3C6D76",
x"8B456D2A",
x"8B846D02",
x"8BF46CF9",
x"8C876D06",
x"8D2B6D21",
x"8DC96D3F",
x"8E506D58",
x"8EB26D69",
x"8EE66D72",
x"8EE76D76",
x"8EC16D7D",
x"8E796D92",
x"8E226DBA",
x"8DCD6DFA",
x"8D8A6E58",
x"8D676ECD",
x"8D6F6F52",
x"8DA56FE1",
x"8E0A7069",
x"8E9470E2",
x"8F397141",
x"8FEC717F",
x"90977197",
x"912B7189",
x"9197715A",
x"91CC710C",
x"91C370A9",
x"917A703A",
x"90F36FC5",
x"90396F55",
x"8F5D6EEF",
x"8E706E99",
x"8D876E59",
x"8CB66E34",
x"8C0D6E2D",
x"8B976E47",
x"8B566E83",
x"8B486EE2",
x"8B636F61",
x"8B9A6FFA",
x"8BDA70A6",
x"8C157157",
x"8C3C71FF",
x"8C45728F",
x"8C2872F4",
x"8BE5731F",
x"8B7F7303",
x"8AFA7296",
x"8A5F71DA",
x"89B270CF",
x"88F96F89",
x"88356E19",
x"876A6C99",
x"86986B26",
x"85BC69D9",
x"84D968CC",
x"83ED680D",
x"82FA67A1",
x"82046786",
x"810E67AE",
x"80206806",
x"7F3E6873",
x"7E7068E1",
x"7DBC6934",
x"7D2B6961",
x"7CC2695E",
x"7C87692E",
x"7C7D68D9",
x"7CA46870",
x"7CFA6806",
x"7D7767AB",
x"7E13676D",
x"7EBB6755",
x"7F626765",
x"7FF36794",
x"805F67D6",
x"8096681D",
x"808D6855",
x"8041686D",
x"7FAC6859",
x"7ED5680E",
x"7DBC678C",
x"7C6666D1",
x"7AD265E2",
x"790064C6",
x"76EF638A",
x"74996231",
x"720060C6",
x"6F285F50",
x"6C1D5DD6",
x"68F55C5D",
x"65CE5AEB",
x"62CB598B",
x"60165843",
x"5DD7571F",
x"5C2E562B",
x"5B34556D",
x"5AF154F1",
x"5B5F54B9",
x"5C6854C9",
x"5DEB551C",
x"5FBE55AE",
x"61B75671",
x"63AB575C",
x"657D585F",
x"6717596A",
x"686F5A71",
x"69875B6A",
x"6A685C4D",
x"6B215D15",
x"6BC25DC2",
x"6C585E56",
x"6CEC5ED7",
x"6D805F4B",
x"6E135FB7",
x"6E9E601F",
x"6F1B6086",
x"6F8560E9",
x"6FD96146",
x"70176198",
x"704A61DC",
x"7077620B",
x"70AD6228",
x"70F76234",
x"715E6235",
x"71E36239",
x"728A624C",
x"734B6279",
x"741A62CC",
x"74EA6349",
x"75AE63EF",
x"765664B5",
x"76DC658B",
x"7737665F",
x"776B6717",
x"777967A1",
x"776D67EC",
x"775167EF",
x"773467A8",
x"77206724",
x"771D666F",
x"7732659E",
x"776064C9",
x"77A46403",
x"77F56359",
x"784962D9",
x"78986281",
x"78D96252",
x"79036243",
x"7911624B",
x"7907625D",
x"78E76277",
x"78BB6290",
x"788A62A8",
x"786262C1",
x"784B62DA",
x"784962FA",
x"78636321",
x"7894634F",
x"78D56381",
x"791A63B4",
x"795563DF",
x"797C63FC",
x"797F6407",
x"795B63FA",
x"790963D8",
x"788E63A1",
x"77F3635C",
x"77426311",
x"768A62CB",
x"75DB6295",
x"753F6276",
x"74C16274",
x"74686291",
x"743162C9",
x"741A6317",
x"741D636F",
x"742E63C2",
x"74476406",
x"745C642A",
x"74666425",
x"746263F2",
x"744C638E",
x"74246300",
x"73EF624F",
x"73AF618A",
x"736D60BF",
x"73316001",
x"73005F5F",
x"72E35EE4",
x"72E05E9A",
x"72FA5E83",
x"73345E9D",
x"738A5EDF",
x"73F95F3E",
x"74765FAB",
x"74FA6015",
x"757A6070",
x"75EF60AF",
x"764C60CC",
x"769060C5",
x"76B8609F",
x"76C56063",
x"76BC601D",
x"76A15FD9",
x"767A5FA7",
x"764B5F8D",
x"76135F94",
x"75D15FB8",
x"757D5FF3",
x"75116037",
x"74836073",
x"73C86095",
x"72D8608B",
x"71AB6048",
x"70445FC1",
x"6E9E5EF3",
x"6CC55DE4",
x"6ABE5C9F",
x"689A5B38",
x"666559C0",
x"64335852",
x"621156FE",
x"601655D9",
x"5E4B54EE",
x"5CC05447",
x"5B7D53E6",
x"5A8A53C4",
x"59E953DE",
x"5997542B",
x"5990549C",
x"59CB5526",
x"5A4155BF",
x"5AE6565D",
x"5BB656F5",
x"5CA45785",
x"5DAE5808",
x"5ED2587E",
x"600C58E7",
x"61565949",
x"62B259A4",
x"64145A01",
x"65765A61",
x"66CC5ACC",
x"680A5B40",
x"69235BBD",
x"6A0F5C3F",
x"6AC95CBF",
x"6B535D32",
x"6BB45D8E",
x"6BF95DC8",
x"6C335DDA",
x"6C725DC1",
x"6CCB5D7B",
x"6D485D17",
x"6DF25CA2",
x"6ECA5C2F",
x"6FC65BD6",
x"70DC5BAF",
x"71F55BCC",
x"72FC5C3B",
x"73DC5CFD",
x"74865E0D",
x"74EC5F59",
x"750A60C6",
x"74E36238",
x"7484638D",
x"73FD64A8",
x"73636572",
x"72CF65DF",
x"725C65F0",
x"721D65B1",
x"72236537",
x"727A649D",
x"73276404",
x"74236389",
x"75656341",
x"76D9633C",
x"786B637F",
x"79FF6404",
x"7B7D64BC",
x"7CCF6594",
x"7DE06675",
x"7EA56746",
x"7F1867F5",
x"7F3A6872",
x"7F1168B1",
x"7EAB68B0",
x"7E1A686F",
x"7D6D67F2",
x"7CB86742",
x"7C09666C",
x"7B686577",
x"7ADC6474",
x"7A636370",
x"79F9627A",
x"799661A1",
x"793060F2",
x"78BB6077",
x"7832603C",
x"77916041",
x"76D86084",
x"760F60FD",
x"753F619B",
x"7479624B",
x"73CB62F6",
x"73426387",
x"72EC63EA",
x"72CE6413",
x"72E563FA",
x"732E63A1",
x"739A6314",
x"7416625F",
x"7490619A",
x"74F060D5",
x"75286024",
x"752B5F95",
x"74F45F31",
x"74865EF8",
x"73EC5EEC",
x"733A5F04",
x"72875F39",
x"71EF5F88",
x"718C5FEA",
x"71736060",
x"71B260E7",
x"724F6181",
x"7342622B",
x"747A62E0",
x"75DC6397",
x"77456441",
x"789364CC",
x"79A1652B",
x"7A53654E",
x"7A98652A",
x"7A6D64BE",
x"79D66414",
x"78EB633B",
x"77C4624C",
x"7681615F",
x"75426090",
x"741D5FED",
x"731E5F83",
x"72445F4F",
x"71825F45",
x"70C25F4D",
x"6FE95F4F",
x"6EDE5F2C",
x"6D895ECF",
x"6BE35E29",
x"69F35D3D",
x"67CE5C15",
x"65975AC9",
x"637C5978",
x"61B15847",
x"60645757",
x"5FBA56C3",
x"5FCE569C",
x"60A656E7",
x"6237579B",
x"646358A8",
x"670759F3",
x"69EF5B5F",
x"6CEC5CD2",
x"6FD25E33",
x"727A5F72",
x"74CE6083",
x"76C16163",
x"784F6217",
x"798462A2",
x"7A6D6310",
x"7B1D6365",
x"7BA363AA",
x"7C1063E2",
x"7C6F6413",
x"7CC9643B",
x"7D23645D",
x"7D7D647C",
x"7DD8649A",
x"7E3164BB",
x"7E8364E2",
x"7EC96510",
x"7F016546",
x"7F226581",
x"7F2A65BF",
x"7F1165F7",
x"7ED66620",
x"7E7C6632",
x"7E036628",
x"7D7665FF",
x"7CDE65B7",
x"7C466556",
x"7BBE64E6",
x"7B4E6473",
x"7AFD6407",
x"7ACF63AF",
x"7AC26373",
x"7ACE6353",
x"7AEA6352",
x"7B0E6369",
x"7B326394",
x"7B4F63CB",
x"7B656409",
x"7B79644B",
x"7B906490",
x"7BB764D9",
x"7BF3652D",
x"7C4E658D",
x"7CC865FD",
x"7D60667D",
x"7E106709",
x"7ECB6799",
x"7F866824",
x"803268A0",
x"80C56901",
x"81356942",
x"817E695E",
x"81A26955",
x"81A56930",
x"819068F5",
x"816D68B4",
x"81496879",
x"812F6855",
x"812A6851",
x"813E6876",
x"817068C8",
x"81BF6947",
x"822869EB",
x"82A36AAB",
x"831F6B7D",
x"83956C51",
x"83F36D17",
x"842F6DBF",
x"84416E3F",
x"84226E89",
x"83D96E96",
x"836A6E63",
x"82E66DF6",
x"825A6D52",
x"81DB6C87",
x"81766BA4",
x"813B6ABA",
x"813169DB",
x"81586917",
x"81AB687F",
x"82206817",
x"82A567E5",
x"832F67E8",
x"83AB6819",
x"8410686F",
x"845568DF",
x"8479695F",
x"847F69E3",
x"846C6A62",
x"844C6AD7",
x"842A6B3D",
x"840D6B90",
x"83FD6BD2",
x"84016BFF",
x"841A6C19",
x"84446C1E",
x"847A6C0F",
x"84B46BE8",
x"84E96BAD",
x"85106B5F",
x"85216B02",
x"85186A9C",
x"84F06A32",
x"84A869D1",
x"8442697A",
x"83BE6937",
x"831B6907",
x"825868E8",
x"816D68D1",
x"804E68B4",
x"7EEC6880",
x"7D356820",
x"7B1A677F",
x"788C668E",
x"75896541",
x"72176393",
x"6E4B618D",
x"6A475F3E",
x"66375CBD",
x"624F5A2C",
x"5EC757AC",
x"5BCC5560",
x"59865367",
x"580D51D8",
x"576850C3",
x"5789502C",
x"5858500F",
x"59AE5061",
x"5B61510C",
x"5D4451FB",
x"5F335319",
x"610F5450",
x"62C5558F",
x"644D56CC",
x"65A457FE",
x"66D65922",
x"67EB5A38",
x"68EF5B3F",
x"69ED5C38",
x"6AF05D21",
x"6BFA5DF6",
x"6D0D5EB1",
x"6E245F4C",
x"6F385FBE",
x"70416000",
x"71316011",
x"71FC5FF0",
x"72965FA2",
x"72F55F35",
x"73165EB5",
x"72F95E35",
x"72A75DC6",
x"72305D7B",
x"71A45D5D",
x"711E5D73",
x"70B25DBB",
x"70765E2B",
x"70765EB7",
x"70B55F4B",
x"712E5FD3",
x"71D3603F",
x"72906083",
x"734F6097",
x"73F96080",
x"747F6045",
x"74D95FF7",
x"750A5FA8",
x"751A5F69",
x"751B5F4D",
x"75245F5D",
x"754B5FA1",
x"759E6017",
x"762D60B8",
x"76F66177",
x"77F5624C",
x"791A6325",
x"7A5263F9",
x"7B8464BF",
x"7C9B6572",
x"7D816610",
x"7E2B669A",
x"7E916714",
x"7EB56783",
x"7EA067E8",
x"7E5D6844",
x"7E006899",
x"7D9D68E5",
x"7D456927",
x"7D06695C",
x"7CEF6983",
x"7D046997",
x"7D48699A",
x"7DB8698A",
x"7E4E696C",
x"7EFD6941",
x"7FBB690D",
x"807968D5",
x"812A68A1",
x"81C36873",
x"82396852",
x"82866842",
x"82A76844",
x"829D685B",
x"826A6881",
x"821A68B5",
x"81B468EF",
x"81436926",
x"80D2694F",
x"806C6962",
x"80146955",
x"7FCF6923",
x"7F9B68C7",
x"7F766844",
x"7F59679B",
x"7F3E66D9",
x"7F206607",
x"7EF76531",
x"7EC46465",
x"7E8463AD",
x"7E386313",
x"7DE0629B",
x"7D7D6249",
x"7D0B621A",
x"7C866207",
x"7BEA620A",
x"7B316217",
x"7A566227",
x"795B6231",
x"78446231",
x"77196224",
x"75EA620B",
x"74C861EC",
x"73C461C9",
x"72EC61A9",
x"7247618E",
x"71D5617A",
x"718C6169",
x"71556152",
x"71176129",
x"70B260E0",
x"700A6069",
x"6F045FB7",
x"6D915EC1",
x"6BB15D84",
x"696C5C0B",
x"66D95A63",
x"641A58A2",
x"615656E6",
x"5EB7554C",
x"5C6253F1",
x"5A7852EB",
x"590C524E",
x"582D521D",
x"57D95256",
x"580A52EB",
x"58B053CA",
x"59B554DA",
x"5B075604",
x"5C8D5730",
x"5E38584F",
x"5FF95953",
x"61C45A3B",
x"63945B05",
x"65695BBB",
x"67415C64",
x"691E5D0A",
x"6B045DB3",
x"6CF55E67",
x"6EED5F27",
x"70EF5FF0",
x"72F560C1",
x"74F96197",
x"76F5626C",
x"78DD633E",
x"7AA8640A",
x"7C4E64D3",
x"7DC6659B",
x"7F0D6662",
x"8020672A",
x"810067F5",
x"81B468BF",
x"82456987",
x"82BC6A47",
x"83276AF6",
x"83916B8D",
x"84036C04",
x"84836C57",
x"85146C7F",
x"85B46C7A",
x"865C6C4E",
x"87046BFD",
x"87A46B90",
x"88326B10",
x"88A86A8F",
x"89046A16",
x"894969B7",
x"897D697D",
x"89AD6976",
x"89E269A7",
x"8A2C6A13",
x"8A946AB5",
x"8B226B89",
x"8BD66C7D",
x"8CAB6D85",
x"8D976E8A",
x"8E886F7F",
x"8F6D7052",
x"903170F9",
x"90C3716E",
x"911471B0",
x"911E71C3",
x"90DC71B0",
x"90567183",
x"8F977145",
x"8EAF7102",
x"8DB270C0",
x"8CB67082",
x"8BCE7048",
x"8B077012",
x"8A6D6FD9",
x"8A076F9D",
x"89D06F58",
x"89C56F0C",
x"89DA6EB7",
x"8A036E5C",
x"8A346E03",
x"8A606DAD",
x"8A806D62",
x"8A8B6D24",
x"8A816CF8",
x"8A626CDC",
x"8A2F6CD2",
x"89ED6CD7",
x"899E6CE8",
x"89456D02",
x"88E46D1E",
x"887A6D3D",
x"88076D57",
x"878D6D69",
x"870A6D75",
x"86866D76",
x"86016D6F",
x"85876D61",
x"85206D4E",
x"84D56D3B",
x"84AF6D2E",
x"84B66D2B",
x"84ED6D3A",
x"85556D5B",
x"85E96D94",
x"86A16DE5",
x"87706E4B",
x"88486EC1",
x"89146F40",
x"89C26FBE",
x"8A427030",
x"8A83708A",
x"8A7C70C3",
x"8A2870D2",
x"898870B7",
x"88A87070",
x"87977006",
x"86696F82",
x"85366EEE",
x"84146E58",
x"83146DCB",
x"82416D4B",
x"81966CD7",
x"81076C65",
x"807D6BE6",
x"7FD36B45",
x"7EE26A6B",
x"7D81693E",
x"7B8E67B2",
x"78F365BE",
x"75A76365",
x"71B560B9",
x"6D3B5DD6",
x"686B5AE1",
x"637F5805",
x"5EBD556A",
x"5A685332",
x"56BD517A",
x"53EE5053",
x"521A4FBD",
x"514B4FB3",
x"517C5025",
x"529250FB",
x"5467521D",
x"56CA5375",
x"598954EB",
x"5C73566E",
x"5F5C57EE",
x"62205960",
x"64A85AB8",
x"66E55BF0",
x"68CF5D00",
x"6A6B5DE0",
x"6BBD5E91",
x"6CCF5F0E",
x"6DAB5F5C",
x"6E5C5F81",
x"6EEB5F88",
x"6F5C5F80",
x"6FB75F74",
x"6FFF5F76",
x"70375F8E",
x"70665FC5",
x"7090601A",
x"70B8608B",
x"70E36110",
x"7119619B",
x"715B6221",
x"71AE6295",
x"721362F0",
x"7287632A",
x"73096344",
x"738E633F",
x"74116323",
x"748762F4",
x"74EA62C2",
x"75326290",
x"755B6268",
x"7565624E",
x"75546242",
x"752E6246",
x"74FD6258",
x"74CE6273",
x"74A76294",
x"749362B9",
x"749662DF",
x"74B16303",
x"74E26327",
x"7525634C",
x"75756374",
x"75CC63A3",
x"762863D8",
x"76866414",
x"76E96455",
x"774F6498",
x"77BE64D8",
x"7835650B",
x"78B4652D",
x"79356537",
x"79B56524",
x"7A2D64F6",
x"7A9764AE",
x"7AF26456",
x"7B3C63F9",
x"7B7C63A3",
x"7BBB6362",
x"7C066344",
x"7C686350",
x"7CE9638D",
x"7D8E63F6",
x"7E566487",
x"7F376535",
x"801E65F0",
x"80F766AA",
x"81AD6752",
x"822A67DF",
x"82626848",
x"824E6889",
x"81EF68A3",
x"8153689A",
x"808C6876",
x"7FAC683E",
x"7ECB67FA",
x"7DF967B1",
x"7D456766",
x"7CB4671B",
x"7C4666D3",
x"7BF7668D",
x"7BBE6645",
x"7B9065FA",
x"7B6665AE",
x"7B39655F",
x"7B076510",
x"7ACF64C5",
x"7A966484",
x"7A5F6452",
x"7A2E6432",
x"7A09642B",
x"79F0643C",
x"79E06466",
x"79D964A1",
x"79D364EA",
x"79C86535",
x"79B16577",
x"798965A8",
x"794E65C1",
x"790365BB",
x"78AD6597",
x"7853655B",
x"7804650D",
x"77CB64B8",
x"77AE6466",
x"77B46420",
x"77D963E8",
x"781163B9",
x"7846638E",
x"785B6353",
x"782D62FA",
x"7796626D",
x"7679619F",
x"74C16087",
x"72655F25",
x"6F725D86",
x"6C005BB9",
x"684159E0",
x"646D5818",
x"60C75684",
x"5D8A553F",
x"5AF55460",
x"592D53F3",
x"584B53F8",
x"58545468",
x"59355533",
x"5AD05642",
x"5CEF577A",
x"5F6258C3",
x"61F05A07",
x"646B5B33",
x"66A95C39",
x"68905D10",
x"6A135DB2",
x"6B315E1E",
x"6BF65E55",
x"6C765E5D",
x"6CCC5E3D",
x"6D135E00",
x"6D655DB1",
x"6DD85D60",
x"6E7C5D1E",
x"6F595CFA",
x"70725D04",
x"71BB5D45",
x"73285DC1",
x"74A55E77",
x"761E5F5D",
x"77796064",
x"78A66177",
x"7991627D",
x"7A376360",
x"7A94640D",
x"7AAE6476",
x"7A906498",
x"7A4C647A",
x"79F26428",
x"799363B8",
x"79416344",
x"790462E3",
x"78E762AB",
x"78ED62AD",
x"791662EC",
x"795F6369",
x"79C96417",
x"7A4F64E5",
x"7AF365BC",
x"7BB46687",
x"7C906735",
x"7D8967B7",
x"7E9D6809",
x"7FC6682D",
x"80FD682D",
x"82396816",
x"836967F7",
x"847F67DF",
x"856967D5",
x"861867DF",
x"868167F7",
x"869E6819",
x"866D6837",
x"85F66845",
x"8545683C",
x"846F681B",
x"838B67E5",
x"82B467A1",
x"82016760",
x"81866737",
x"81526732",
x"81696760",
x"81C867C5",
x"8263685F",
x"83286920",
x"83FF69F7",
x"84CF6ACF",
x"85806B93",
x"86006C30",
x"86456C9D",
x"864B6CD8",
x"86176CE6",
x"85B66CD7",
x"853B6CB7",
x"84BA6C9C",
x"84466C90",
x"83F46C9D",
x"83D06CC4",
x"83E36D00",
x"842F6D48",
x"84AC6D8F",
x"85526DC8",
x"86106DEC",
x"86CF6DF5",
x"877E6DE2",
x"880B6DBB",
x"88636D85",
x"887E6D4B",
x"885A6D14",
x"88006CE9",
x"877D6CCD",
x"86EA6CC2",
x"86636CCD",
x"86076CE9",
x"85F06D1C",
x"86356D65",
x"86DF6DC7",
x"87EC6E43",
x"89526ED7",
x"8AF96F80",
x"8CC1703A",
x"8E8870F8",
x"903171AF",
x"919B724E",
x"92B472C8",
x"936F7310",
x"93C5731F",
x"93B672EC",
x"9343727C",
x"926C71CD",
x"912B70E4",
x"8F7C6FC7",
x"8D556E78",
x"8AAC6CF9",
x"877D6B4E",
x"83CC697A",
x"7FA76780",
x"7B276569",
x"76736341",
x"71BE6117",
x"6D3E5F01",
x"69275D15",
x"65AD5B6A",
x"62F15A12",
x"6109591C",
x"5FFA588E",
x"5FB85863",
x"6027588F",
x"61245901",
x"628359A1",
x"641C5A53",
x"65C95B04",
x"67705BA1",
x"69005C21",
x"6A735C82",
x"6BCB5CCD",
x"6D105D0D",
x"6E4C5D4F",
x"6F8A5DA5",
x"70CF5E1A",
x"721A5EB3",
x"73665F70",
x"74A8604B",
x"75D66137",
x"76E56224",
x"77CB6304",
x"788A63CF",
x"7928647F",
x"79B16511",
x"7A34658E",
x"7AC16600",
x"7B656670",
x"7C2466E5",
x"7CFC6760",
x"7DD967E0",
x"7EA86858",
x"7F4968BA",
x"7F9E68F3",
x"7F9068F5",
x"7F0D68B4",
x"7E13682D",
x"7CAF6766",
x"7AFD666D",
x"79216558",
x"7745643F",
x"7597633E",
x"74396268",
x"734761CE",
x"72CC6179",
x"72C76168",
x"73286197",
x"73D961FA",
x"74BA6289",
x"75AD6332",
x"769963F0",
x"776964B8",
x"78116584",
x"7890664F",
x"78E76714",
x"792567D1",
x"7955687C",
x"79806911",
x"79B26989",
x"79F269E1",
x"7A3F6A13",
x"7A9D6A21",
x"7B036A11",
x"7B6F69EC",
x"7BDB69BC",
x"7C41698E",
x"7C9E696F",
x"7CF36968",
x"7D3F697F",
x"7D8369B7",
x"7DBC6A0F",
x"7DED6A7C",
x"7E136AF5",
x"7E276B6D",
x"7E2A6BD7",
x"7E176C24",
x"7DF26C4E",
x"7DBC6C4F",
x"7D836C28",
x"7D536BE1",
x"7D446B80",
x"7D656B17",
x"7DCC6AB1",
x"7E846A5C",
x"7F946A21",
x"80F06A06",
x"82866A06",
x"84356A1C",
x"85D26A3B",
x"87326A56",
x"882D6A61",
x"889F6A4E",
x"88796A1A",
x"87B969C7",
x"86746958",
x"84CF68DE",
x"82FC6862",
x"812F67F7",
x"7FA167A8",
x"7E7F677D",
x"7DE26777",
x"7DD66793",
x"7E4F67C9",
x"7F31680E",
x"80516856",
x"81806897",
x"829068CB",
x"835C68EF",
x"83CE6906",
x"83DD6913",
x"8395691D",
x"830B6928",
x"82606937",
x"81B26948",
x"811A6955",
x"80A46952",
x"80526934",
x"801068EB",
x"7FBF6869",
x"7F3B67A7",
x"7E5B66A1",
x"7CFD6556",
x"7B0E63D2",
x"788A6221",
x"75846058",
x"72235E88",
x"6E995CCD",
x"6B245B3B",
x"680559E1",
x"657058D0",
x"6392580F",
x"627F579F",
x"623B577E",
x"62B657A2",
x"63CC5801",
x"6557588B",
x"67255932",
x"690F59E9",
x"6AF05AA2",
x"6CB35B57",
x"6E4A5C04",
x"6FBA5CA8",
x"710A5D48",
x"724C5DE7",
x"73905E91",
x"74E55F4C",
x"7652601F",
x"77DB6111",
x"7979621F",
x"7B216348",
x"7CC46483",
x"7E5365C4",
x"7FBF66FA",
x"80FC681A",
x"82036913",
x"82D369D9",
x"83726A66",
x"83E56AB5",
x"84376ACB",
x"84766AAE",
x"84AE6A6B",
x"84E96A10",
x"853169B0",
x"858D6958",
x"86036919",
x"869468FD",
x"8742690D",
x"880B694C",
x"88EF69BC",
x"89E76A59",
x"8AF16B1E",
x"8C066C03",
x"8D1B6CFD",
x"8E2E6E03",
x"8F386F0A",
x"90327008",
x"912170F6",
x"920471CE",
x"92E4728F",
x"93CB7339",
x"94C173CD",
x"95D07452",
x"96FD74CB",
x"9848753D",
x"99A975A6",
x"9B117603",
x"9C6C7650",
x"9D9F7682",
x"9E95768D",
x"9F35766A",
x"9F6E760F",
x"9F3E757C",
x"9EA574B9",
x"9DB673D1",
x"9C8D72D8",
x"9B4671E6",
x"9A077114",
x"98F17075",
x"98217017",
x"97A57000",
x"97817027",
x"97AC707F",
x"981470EF",
x"9898715B",
x"991871AB",
x"997371CB",
x"998E71AF",
x"99577157",
x"98C870CD",
x"97EA7026",
x"96D26F7C",
x"959A6EE8",
x"94666E80",
x"93566E55",
x"92836E6B",
x"91FD6EBA",
x"91C56F31",
x"91C96FB7",
x"91F3702E",
x"9218707A",
x"92157085",
x"91C3703B",
x"91076F9A",
x"8FD86EAB",
x"8E396D7F",
x"8C466C31",
x"8A286AE2",
x"881069AE",
x"863268B4",
x"84BE6809",
x"83D567B5",
x"838767BE",
x"83D06814",
x"849568A6",
x"85AF6959",
x"86EA6A13",
x"88116AB8",
x"88F76B32",
x"897D6B78",
x"89906B82",
x"89356B57",
x"887E6B02",
x"878A6A94",
x"86796A21",
x"856A69B5",
x"8470695C",
x"83916916",
x"82BF68DB",
x"81E3689B",
x"80D66842",
x"7F7367BA",
x"7D9A66EC",
x"7B3465CC",
x"78426453",
x"74D66289",
x"71166077",
x"6D3A5E3D",
x"697D5BF8",
x"662359CD",
x"635F57DD",
x"615B5644",
x"6029551B",
x"5FC55468",
x"601C5430",
x"61095467",
x"625B54FB",
x"63E655D3",
x"657D56D6",
x"670057E7",
x"685E58F1",
x"698D59E1",
x"6A945AAC",
x"6B805B4F",
x"6C625BC9",
x"6D485C24",
x"6E3B5C69",
x"6F415CA8",
x"70515CEC",
x"71655D3C",
x"726D5DA2",
x"735E5E1F",
x"742A5EB1",
x"74CB5F4F",
x"75415FF6",
x"75936098",
x"75C96131",
x"75F361B7",
x"761E6225",
x"7658627E",
x"76A762C1",
x"770E62F0",
x"778D6313",
x"781B632D",
x"78B26341",
x"79476353",
x"79CE6366",
x"7A44637A",
x"7AA3638E",
x"7AEC63A3",
x"7B2163B8",
x"7B4863CE",
x"7B6663E3",
x"7B8163FC",
x"7BA16417",
x"7BC96437",
x"7BFF645A",
x"7C426486",
x"7C9964BA",
x"7D0464F9",
x"7D8A6546",
x"7E2B65A5",
x"7EE9661A",
x"7FC866A7",
x"80C5674B",
x"81DC6806",
x"830968D2",
x"844269AB",
x"857D6A87",
x"86B26B5E",
x"87D96C23",
x"88EA6CD2",
x"89E66D66",
x"8ACC6DE1",
x"8BA16E45",
x"8C6C6E9A",
x"8D326EE8",
x"8DF66F35",
x"8EB96F89",
x"8F776FE4",
x"90277043",
x"90B8709F",
x"911D70EC",
x"9142711F",
x"911A7126",
x"909A70F8",
x"8FBB708F",
x"8E836FE8",
x"8CF96F0A",
x"8B316DFF",
x"893F6CD7",
x"873E6BA7",
x"85466A83",
x"8373697F",
x"81D568AA",
x"807E680D",
x"7F7567AD",
x"7EBA6787",
x"7E456790",
x"7E0B67BE",
x"7DFD67FC",
x"7E0B683E",
x"7E246872",
x"7E3C6890",
x"7E4F6891",
x"7E5C687A",
x"7E69684F",
x"7E83681E",
x"7EB867F5",
x"7F1767E2",
x"7FAA67F0",
x"80766826",
x"81746883",
x"829B6900",
x"83D3698E",
x"85016A1E",
x"860B6A9C",
x"86D66AF5",
x"87516B1A",
x"87706B07",
x"87376ABD",
x"86B46A42",
x"85F769A7",
x"851B68FA",
x"8431684E",
x"834567AE",
x"82596723",
x"816566AD",
x"80526642",
x"7F0A65DB",
x"7D706568",
x"7B7664DA",
x"7916642B",
x"765C635A",
x"736A626F",
x"70726179",
x"6DAE6090",
x"6B615FCB",
x"69C55F46",
x"69075F17",
x"69445F49",
x"6A7D5FE2",
x"6CA060DC",
x"6F866228",
x"72FC63B4",
x"76C96569",
x"7AB96732",
x"7EA068FD",
x"825D6ABE",
x"85E56C70",
x"89356E10",
x"8C566FA4",
x"8F5A712E",
x"925672B6",
x"9559743D",
x"986E75C3",
x"9BA27746",
x"9EF178C0",
x"A25C7A2D",
x"A5DA7B88",
x"A9637CCA",
x"ACE87DF2",
x"B05D7EFE",
x"B3B57FF0",
x"B6DA80C6",
x"B9BD8185",
x"BC4C822D",
x"BE7782C0",
x"C033833F",
x"C17B83AB",
x"C2538401",
x"C2C48446",
x"C2E18478",
x"C2C3849B",
x"C28284AD",
x"C23984B6",
x"C1F884B6",
x"C1D084B1",
x"C1C484A9",
x"C1D384A2",
x"C1F484A3",
x"C21984AF",
x"C23A84CD",
x"C24E8501",
x"C2518552",
x"C24685C0",
x"C235864D",
x"C22886F1",
x"C22C87A5",
x"C250885F",
x"C298890E",
x"C30889A8",
x"C3998A1D",
x"C43D8A64",
x"C4E38A79",
x"C56F8A56",
x"C5CB8A03",
x"C5E18983",
x"C59B88E2",
x"C4EB8827",
x"C3CE875C",
x"C249868A",
x"C06785B5",
x"BE3F84E6",
x"BBED841E",
x"B9948363",
x"B75482BB",
x"B554822C",
x"B3B281C2",
x"B2828185",
x"B1D4817D",
x"B1AC81AF",
x"B1FE821C",
x"B2B982C2",
x"B3C28394",
x"B4F78481",
x"B6388577",
x"B764865D",
x"B8638721",
x"B91E87AE",
x"B98F87F7",
x"B9B587F9",
x"B99487B3",
x"B9398732",
x"B8AD8683",
x"B7FE85B8",
x"B72D84E3",
x"B63A840F",
x"B51F834A",
x"B3D08294",
x"B24281E7",
x"B069813B",
x"AE3C8081",
x"ABC27FAD",
x"A8FE7EB5",
x"A6087D91",
x"A2F87C44",
x"9FF37ADA",
x"9D1A7962",
x"9A8D77F2",
x"986776A5",
x"96BC758D",
x"959474BD",
x"94E47439",
x"94A173FF",
x"94AC7400",
x"94E77426",
x"952B7454",
x"9556746E",
x"95487457",
x"94EC73FC",
x"94327354",
x"9318725F",
x"91A5712A",
x"8FE96FC8",
x"8DF66E4E",
x"8BDF6CD2",
x"89B76B68",
x"87886A1A",
x"855668E9",
x"831B67CC",
x"80C966BA",
x"7E4E659B",
x"7B966460",
x"789062FD",
x"75376168",
x"718C5FA4",
x"6DA15DBB",
x"69945BBD",
x"658F59C7",
x"61BD57EE",
x"5E52564F",
x"5B7954FA",
x"595253FF",
x"57F35367",
x"57615330",
x"578D5354",
x"586253C7",
x"59BD5477",
x"5B755554",
x"5D61564F",
x"5F5F5753",
x"614F5856",
x"631C594D",
x"64B85A30",
x"661E5AF8",
x"67515BA5",
x"68545C35",
x"69305CAB",
x"69ED5D0A",
x"6A935D57",
x"6B285D97",
x"6BB25DCF",
x"6C335E04",
x"6CAB5E38",
x"6D1E5E6E",
x"6D8C5EA5",
x"6DF25ED9",
x"6E525F08",
x"6EAD5F2F",
x"6F025F48",
x"6F525F52",
x"6FA05F4B",
x"6FEC5F35",
x"703C5F12",
x"70945EEA",
x"70F55EC1",
x"71625E9B",
x"71DB5E7D",
x"725D5E69",
x"72E35E5F",
x"73685E5C",
x"73DF5E59",
x"74445E55",
x"748D5E49",
x"74B55E33",
x"74BD5E14",
x"74A45DEE",
x"74705DC8",
x"74275DA8",
x"73D35D98",
x"737A5D9C",
x"73245DB9",
x"72D25DEE",
x"72895E36",
x"72455E87",
x"72075ED6",
x"71CF5F18",
x"719D5F46",
x"71725F5A",
x"71565F55",
x"71515F3F",
x"716B5F22",
x"71AA5F0E",
x"72135F12",
x"72A85F3B",
x"73635F8E",
x"743B600D",
x"752060B2",
x"75FD616F",
x"76C26231",
x"775B62E6",
x"77BA637A",
x"77D663E2",
x"77AE6413",
x"7748640E",
x"76B163D9",
x"75FA6383",
x"7538631A",
x"748262AE",
x"73E96250",
x"737C620B",
x"734461E8",
x"734161E6",
x"736F6204",
x"73C26239",
x"742D627C",
x"749D62BF",
x"750262F9",
x"754C631F",
x"7575632A",
x"75756313",
x"754C62DA",
x"75026283",
x"749E6211",
x"742D618D",
x"73BA60FE",
x"734E6072",
x"72EF5FEE",
x"72A15F7E",
x"72635F22",
x"72325EDF",
x"72065EB1",
x"71D85E92",
x"71A15E7D",
x"715C5E6A",
x"71045E52",
x"709A5E33",
x"701E5E0E",
x"6F965DE4",
x"6F035DBF",
x"6E6D5DA5",
x"6DDB5D9F",
x"6D4B5DB1",
x"6CC25DDD",
x"6C415E1E",
x"6BC25E6A",
x"6B425EB1",
x"6ABB5EE3",
x"6A265EED",
x"697B5EBF",
x"68B45E4F",
x"67D15D95",
x"66D15C9A",
x"65BA5B63",
x"64935A07",
x"6366589A",
x"62425735",
x"613355F1",
x"604454E6",
x"5F7D5423",
x"5EE553B6",
x"5E7C53A1",
x"5E4353E1",
x"5E315470",
x"5E48553D",
x"5E82563C",
x"5EDC5759",
x"5F5B5882",
x"600059AB",
x"60D25AC5",
x"61D85BC9",
x"63135CB1",
x"64865D7A",
x"66305E24",
x"68065EAE",
x"6A025F1E",
x"6C145F76",
x"6E335FBE",
x"704F5FFC",
x"72616039",
x"74606080",
x"764A60DA",
x"781B6155",
x"79D661F7",
x"7B7A62C8",
x"7D0963C5",
x"7E7D64E8",
x"7FD56624",
x"81086763",
x"8214688E",
x"82F0698D",
x"839A6A47",
x"84106AAB",
x"84526AB4",
x"84656A63",
x"844E69C5",
x"841568F2",
x"83C26803",
x"835A6716",
x"82E66642",
x"826A659B",
x"81EA652A",
x"817064ED",
x"80FD64DF",
x"809B64EC",
x"804F6507",
x"801E651E",
x"800D6527",
x"801B651D",
x"80486501",
x"808C64DC",
x"80DF64BA",
x"813864A7",
x"818B64AF",
x"81D064DA",
x"81FE652A",
x"8214659B",
x"820E6625",
x"81F066BC",
x"81BE6755",
x"817C67E2",
x"812F685B",
x"80E268BA",
x"809768FA",
x"8056691E",
x"80276928",
x"8013691D",
x"80216903",
x"805D68DE",
x"80CC68B4",
x"8173688A",
x"82506865",
x"835F6849",
x"8491683E",
x"85D56845",
x"87166866",
x"883E68A6",
x"893B6907",
x"89FE698C",
x"8A866A32",
x"8AD26AF5",
x"8AF06BCA",
x"8AF16CA6",
x"8AE76D79",
x"8AE36E34",
x"8AF36ECA",
x"8B1A6F2B",
x"8B566F52",
x"8B9D6F3B",
x"8BDD6EE9",
x"8C096E65",
x"8C106DBA",
x"8BE96CF9",
x"8B956C33",
x"8B1B6B76",
x"8A8A6AD1",
x"89F66A4C",
x"897369EF",
x"891569BA",
x"88ED69AD",
x"890169C4",
x"895069FA",
x"89D26A4B",
x"8A776AB0",
x"8B2F6B23",
x"8BE66BA0",
x"8C8B6C20",
x"8D126C9E",
x"8D766D17",
x"8DB56D83",
x"8DD56DE1",
x"8DDD6E2B",
x"8DD66E62",
x"8DC66E83",
x"8DAE6E8D",
x"8D866E80",
x"8D416E58",
x"8CC86E0F",
x"8BFD6D9C",
x"8AC16CF2",
x"88F46C06",
x"867C6AC9",
x"83466932",
x"7F52673C",
x"7AAB64E9",
x"75706241",
x"6FD25F5A",
x"6A0D5C4F",
x"64635943",
x"5F1D565A",
x"5A7B53BA",
x"56B15185",
x"53E94FD3",
x"52344EB3",
x"518F4E2A",
x"51E64E33",
x"53174EBC",
x"54F24FAD",
x"574550EA",
x"59DE5257",
x"5C9053D6",
x"5F3A554E",
x"61C056B0",
x"641357EE",
x"662B5902",
x"680759EE",
x"69AB5AB5",
x"6B195B5D",
x"6C555BF0",
x"6D635C76",
x"6E455CF7",
x"6EFD5D7A",
x"6F905E03",
x"70015E95",
x"70595F32",
x"709E5FD9",
x"70DB6088",
x"7116613B",
x"715861ED",
x"71A36295",
x"71F9632F",
x"725663AF",
x"72B76410",
x"73166448",
x"736C6458",
x"73B5643B",
x"73F363F7",
x"74246391",
x"744C6315",
x"74736290",
x"749E620D",
x"74D2619B",
x"75146146",
x"75636114",
x"75BF610A",
x"76236125",
x"76876162",
x"76E961B7",
x"77416218",
x"778E627A",
x"77D162D5",
x"780D631D",
x"784C634F",
x"7897636C",
x"78FA6374",
x"797F6372",
x"7A2A6369",
x"7AFD6368",
x"7BF46374",
x"7D036397",
x"7E1A63D5",
x"7F25642F",
x"800D64A3",
x"80C1652B",
x"812F65C1",
x"81536660",
x"812E66FF",
x"80CE679B",
x"80466831",
x"7FB568C1",
x"7F3E694C",
x"7F0069D6",
x"7F166A63",
x"7F966AF3",
x"80866B86",
x"81E06C1D",
x"83936CB1",
x"85806D3E",
x"87816DBB",
x"89706E23",
x"8B286E6E",
x"8C876E99",
x"8D796EA1",
x"8DF36E88",
x"8DF66E4E",
x"8D916DFA",
x"8CD56D96",
x"8BDA6D26",
x"8ABB6CB3",
x"898B6C44",
x"885A6BE2",
x"87376B92",
x"86216B54",
x"851E6B2D",
x"842C6B19",
x"834E6B14",
x"82816B17",
x"81CF6B1D",
x"813F6B1D",
x"80DC6B10",
x"80AE6AF0",
x"80B96ABF",
x"81036A7A",
x"81816A2A",
x"822B69D5",
x"82EC6984",
x"83AF6942",
x"84636919",
x"84F4690A",
x"8559691B",
x"8593694B",
x"85A56994",
x"85A069ED",
x"85916A4E",
x"85876AA7",
x"858A6AEF",
x"85986B19",
x"85A46B1A",
x"85956AE9",
x"854E6A80",
x"84AA69D9",
x"838B68F5",
x"81DF67D3",
x"7F9D667D",
x"7CD564FD",
x"79A56366",
x"764161C9",
x"72E0603F",
x"6FC65EDD",
x"6D2D5DBB",
x"6B455CE4",
x"6A2E5C69",
x"69F05C46",
x"6A835C7B",
x"6BC95CFA",
x"6D975DB2",
x"6FBE5E92",
x"720D5F8B",
x"745B608B",
x"7689618D",
x"78896289",
x"7A536381",
x"7BF3647A",
x"7D776575",
x"7EF16675",
x"80736779",
x"82096881",
x"83B76986",
x"857B6A83",
x"87516B72",
x"89296C4F",
x"8AFA6D1D",
x"8CB96DDE",
x"8E606E99",
x"8FEC6F58",
x"915F7021",
x"92BF70FC",
x"941171E8",
x"955A72E1",
x"969D73DB",
x"97D374CB",
x"98FD75A2",
x"9A0E7652",
x"9B0176D2",
x"9BCF7720",
x"9C78773C",
x"9D01772F",
x"9D717706",
x"9DD976D0",
x"9E457699",
x"9EC87672",
x"9F6C7660",
x"A0357667",
x"A1257686",
x"A23076BC",
x"A34B76FF",
x"A45F774A",
x"A55A7799",
x"A62E77E7",
x"A6CF7834",
x"A73A7882",
x"A77778D3",
x"A792792C",
x"A7A17990",
x"A7B67A03",
x"A7E97A89",
x"A8477B22",
x"A8DF7BCC",
x"A9AB7C81",
x"AAA37D3D",
x"ABB97DF8",
x"ACD27EA9",
x"ADD27F42",
x"AEA67FBD",
x"AF3A8012",
x"AF81803D",
x"AF7D803C",
x"AF368015",
x"AEC07FD3",
x"AE357F82",
x"ADAE7F36",
x"AD467EFE",
x"AD117EE8",
x"AD157EFE",
x"AD567F46",
x"ADC67FBD",
x"AE548057",
x"AEE98107",
x"AF6981B6",
x"AFC08256",
x"AFE382D1",
x"AFCA8321",
x"AF78833B",
x"AEF88321",
x"AE5A82D7",
x"ADAB826A",
x"ACF881E3",
x"AC45814C",
x"AB8F80AF",
x"AACF800F",
x"A9F47F6E",
x"A8EE7EC9",
x"A7AE7E18",
x"A6267D57",
x"A4597C81",
x"A24D7B92",
x"A0147A8C",
x"9DC97975",
x"9B8D7856",
x"9983773D",
x"97CC7639",
x"96807558",
x"95B174A6",
x"9562742F",
x"958673F2",
x"960873F2",
x"96CB7423",
x"97A5747C",
x"987374EC",
x"99127562",
x"996A75CE",
x"996F7623",
x"9924765B",
x"98957671",
x"97DF7668",
x"971B7644",
x"9664760C",
x"95CF75C6",
x"955D7574",
x"95047512",
x"94A47499",
x"941173FE",
x"931B7330",
x"918B721F",
x"8F3970C0",
x"8C0D6F0A",
x"88066CFF",
x"833E6AA8",
x"7DE5681B",
x"78456573",
x"72B062CE",
x"6D7C604F",
x"68F75E15",
x"65635C3D",
x"62E85AD9",
x"619159F3",
x"61595988",
x"621D5992",
x"63B059FE",
x"65D25AB9",
x"684C5BA5",
x"6AE25CAC",
x"6D655DB3",
x"6FAD5EA7",
x"71A45F78",
x"733F601F",
x"747F609D",
x"756D60F2",
x"761D612E",
x"76A5615F",
x"771D6195",
x"779A61E4",
x"78306256",
x"78EC62F3",
x"79D363BC",
x"7AE564AA",
x"7C1365B1",
x"7D4C66BF",
x"7E7F67C4",
x"7F9168AD",
x"806F696C",
x"810469F9",
x"814B6A4F",
x"813F6A75",
x"80E96A6F",
x"80536A48",
x"7F946A0C",
x"7EBE69C4",
x"7DE66976",
x"7D206927",
x"7C7768D6",
x"7BF46884",
x"7B9A682D",
x"7B6367CE",
x"7B4C6769",
x"7B4B66FF",
x"7B596696",
x"7B6D6634",
x"7B8465E3",
x"7B9D65AA",
x"7BB76591",
x"7BD5659B",
x"7BFF65CC",
x"7C376623",
x"7C83669A",
x"7CE9672D",
x"7D6967CF",
x"7E016877",
x"7EB0691B",
x"7F6A69B0",
x"80286A27",
x"80D96A7A",
x"816F6AA3",
x"81DC6A9C",
x"82146A66",
x"820E6A06",
x"81C66984",
x"813E68EC",
x"807D6846",
x"7F9167A4",
x"7E8D670D",
x"7D816689",
x"7C84661E",
x"7BA565CB",
x"7AF2658E",
x"7A72655F",
x"7A25653B",
x"7A0C6518",
x"7A1764F4",
x"7A4164CE",
x"7A7764A5",
x"7AB1647F",
x"7AE2645D",
x"7AFE6445",
x"7B046439",
x"7AED6437",
x"7AB96439",
x"7A69643C",
x"79FF6432",
x"797F6415",
x"78EB63DF",
x"784B638A",
x"77A56317",
x"7700628E",
x"766361F7",
x"75D86160",
x"756260D6",
x"75066067",
x"74C7601B",
x"74A35FFC",
x"74946007",
x"7496603B",
x"749B6090",
x"749B60FA",
x"7490616D",
x"746F61DD",
x"7435623C",
x"73E36281",
x"737962A2",
x"72FA629A",
x"726B6264",
x"71D16201",
x"712D6174",
x"708160C3",
x"6FCE5FF6",
x"6F105F1A",
x"6E475E39",
x"6D6F5D64",
x"6C8A5CA7",
x"6B975C0A",
x"6A9A5B92",
x"69965B3F",
x"688D5B0B",
x"67865AEB",
x"66835AD3",
x"65865AAF",
x"64905A74",
x"63A15A18",
x"62BA5995",
x"61DE58F3",
x"610C5836",
x"604C5774",
x"5FA656BF",
x"5F1E562B",
x"5EBE55C9",
x"5E8D55A5",
x"5E9055C6",
x"5EC75628",
x"5F3356C2",
x"5FCE5784",
x"6090585D",
x"61735939",
x"626D5A08",
x"63785AC0",
x"648C5B59",
x"65A65BD0",
x"66C25C29",
x"67E35C6D",
x"69055CA1",
x"6A275CD0",
x"6B485D01",
x"6C635D3B",
x"6D755D80",
x"6E735DD2",
x"6F5C5E32",
x"70275E9D",
x"70D15F0D",
x"71565F7D",
x"71B85FE7",
x"71F96045",
x"721D608E",
x"723060BE",
x"723560D0",
x"723D60C6",
x"724F60A1",
x"7277606A",
x"72C1602E",
x"73325FF9",
x"73D25FD9",
x"74A05FDF",
x"759B6010",
x"76BC6073",
x"77F96104",
x"794261BB",
x"7A8D6289",
x"7BC6635D",
x"7CE56425",
x"7DDF64D0",
x"7EB16552",
x"7F5C65A5",
x"7FE365CC",
x"805265CE",
x"80B265BB",
x"810E65A3",
x"816F659A",
x"81DB65AF",
x"825265F3",
x"82D5666A",
x"835F6717",
x"83E767F0",
x"846968EB",
x"84DC69F5",
x"853C6AFC",
x"858A6BED",
x"85C66CBD",
x"85F66D5C",
x"86206DCA",
x"864E6E0A",
x"86886E26",
x"86DB6E2D",
x"87486E2D",
x"87D86E35",
x"88886E55",
x"89586E90",
x"8A3F6EE5",
x"8B346F4D",
x"8C276FBA",
x"8D0D701F",
x"8DD6706B",
x"8E777094",
x"8EE97096",
x"8F247073",
x"8F297034",
x"8EFE6FEC",
x"8EAC6FAA",
x"8E3B6F82",
x"8DB66F7E",
x"8D2A6FA6",
x"8C9D6FF5",
x"8C11705F",
x"8B8B70D2",
x"8B097137",
x"8A837175",
x"89F67179",
x"895C7134",
x"88B470A3",
x"87FA6FCA",
x"87346EB4",
x"86676D76",
x"859E6C2A",
x"84E26AE6",
x"843C69C4",
x"83B768D6",
x"8356682A",
x"831A67C6",
x"82FC67AA",
x"82F467CF",
x"82F46827",
x"82ED68A4",
x"82D06932",
x"829369BE",
x"822A6A37",
x"81936A8D",
x"80D16AB5",
x"7FE96AA7",
x"7EE76A61",
x"7DD569E3",
x"7CBC6937",
x"7BA76866",
x"7A97677C",
x"798A6686",
x"787D6590",
x"776564A4",
x"763863C8",
x"74F26301",
x"738D6252",
x"720D61B7",
x"7079612D",
x"6EE360AF",
x"6D5F603E",
x"6C045FD8",
x"6AEB5F7C",
x"6A285F2F",
x"69CC5EF7",
x"69DF5ED7",
x"6A5E5ED9",
x"6B415EFD",
x"6C7A5F45",
x"6DF65FB1",
x"6F9B603C",
x"715860DF",
x"73176193",
x"74CE624E",
x"76706309",
x"780063BF",
x"797A646C",
x"7AE5650D",
x"7C4165A3",
x"7D93662D",
x"7ED866AE",
x"800E6725",
x"812F6794",
x"823467F9",
x"83146852",
x"83C968A1",
x"845268E5",
x"84AF691E",
x"84E66952",
x"85006984",
x"850769BB",
x"850A69FA",
x"85106A48",
x"85226AA3",
x"85456B0A",
x"85766B75",
x"85B46BDC",
x"85F66C34",
x"86326C70",
x"86636C89",
x"86816C76",
x"868A6C37",
x"867E6BD1",
x"86656B4F",
x"86456AC2",
x"862E6A3A",
x"862C69CB",
x"864F6984",
x"86A06972",
x"8728699A",
x"87EC69FA",
x"88E66A8D",
x"8A0E6B45",
x"8B596C16",
x"8CB66CF0",
x"8E146DC7",
x"8F606E8F",
x"908E6F44",
x"91916FE2",
x"92647069",
x"930570DA",
x"93777133",
x"93C07174",
x"93E77197",
x"93F9719D",
x"93F97182",
x"93F07141",
x"93E170E1",
x"93D07065",
x"93B96FD7",
x"939E6F45",
x"93796EBF",
x"93466E4F",
x"93056E02",
x"92B66DD8",
x"92556DCF",
x"91E26DDF",
x"915F6DFA",
x"90CC6E0F",
x"902E6E0C",
x"8F846DE6",
x"8ED06D97",
x"8E176D1D",
x"8D566C80",
x"8C936BCC",
x"8BC86B13",
x"8AF96A65",
x"8A2569CF",
x"8949695F",
x"88676919",
x"877C68FA",
x"868A68FC",
x"858E6911",
x"848D692B",
x"8383693A",
x"8277692E",
x"816968FC",
x"805F68A0",
x"7F5D6819",
x"7E6C676D",
x"7D9466A8",
x"7CDE65DB",
x"7C526514",
x"7BF66468",
x"7BCE63E5",
x"7BD66397",
x"7C096381",
x"7C5863A1",
x"7CB463ED",
x"7D046456",
x"7D3764C9",
x"7D386534",
x"7CFC6581",
x"7C7D65A4",
x"7BC26593",
x"7AD8654C",
x"79D164D2",
x"78C5642F",
x"77C6636D",
x"76E8629A",
x"762A61BC",
x"758960E0",
x"74F26004",
x"74475F2B",
x"73665E4D",
x"72305D69",
x"70865C77",
x"6E565B74",
x"6BA05A60",
x"68735942",
x"64EC581E",
x"613A5702",
x"5D9255FA",
x"5A275514",
x"57305459",
x"54D553D3",
x"53335388",
x"52555378",
x"523953A2",
x"52CD53FF",
x"53F55487",
x"55925532",
x"577C55F4",
x"599256C3",
x"5BB75797",
x"5DD15863",
x"5FCC5922",
x"61A059D2",
x"63415A6B",
x"64AB5AF4",
x"65E15B6A",
x"66DF5BD6",
x"67AD5C3D",
x"684C5CA4",
x"68C55D11",
x"691E5D84",
x"69615E00",
x"69945E7C",
x"69C15EF1",
x"69EB5F56",
x"6A145F9F",
x"6A3F5FC2",
x"6A665FB9",
x"6A865F83",
x"6A975F21",
x"6A965E9D",
x"6A7D5E04",
x"6A4C5D64",
x"6A075CCD",
x"69B45C4F",
x"695B5BF3",
x"69055BBB",
x"68BE5BA9",
x"688F5BB6",
x"687A5BDA",
x"68875C07",
x"68B45C31",
x"68FD5C4C",
x"695F5C55",
x"69D15C48",
x"6A515C26",
x"6AD85BF8",
x"6B655BC9",
x"6BF85BA4",
x"6C905B98",
x"6D335BAF",
x"6DDE5BF3",
x"6E975C66",
x"6F5B5D07",
x"70285DCF",
x"70F95EAF",
x"71C55F98",
x"72836077",
x"73286139",
x"73AB61CE",
x"74026228",
x"74276242",
x"7419621F",
x"73DB61C6",
x"73756142",
x"72F060A7",
x"725B6004",
x"71C25F6C",
x"71345EEC",
x"70BB5E90",
x"705F5E5A",
x"70215E4D",
x"70005E63",
x"6FF65E94",
x"6FFC5ED6",
x"700A5F22",
x"70195F70",
x"70245FBE",
x"702A6007",
x"702A604D",
x"70276091",
x"702360D5",
x"70216117",
x"70236156",
x"70246190",
x"702061BB",
x"701161D3",
x"6FF361CF",
x"6FBB61A9",
x"6F68615D",
x"6EF560E9",
x"6E63604F",
x"6DB75F95",
x"6CF55EC6",
x"6C235DED",
x"6B485D15",
x"6A695C4C",
x"698D5B9A",
x"68BA5B07",
x"67F35A97",
x"673F5A4A",
x"66A95A1F",
x"66345A14",
x"65EC5A21",
x"65D75A42",
x"65F65A71",
x"664A5AAC",
x"66C75AF0",
x"67645B38",
x"68075B81",
x"689D5BC8",
x"690C5C08",
x"693C5C3D",
x"69205C61",
x"68AE5C6E",
x"67EE5C60",
x"66EB5C36",
x"65BE5BF1",
x"64835B92",
x"63585B21",
x"62565AA4",
x"61905A21",
x"610C59A2",
x"60C2592B",
x"60A658BD",
x"6099585C",
x"60805804",
x"603D57AF",
x"5FBB575D",
x"5EEF570A",
x"5DDB56B5",
x"5C905661",
x"5B2B5616",
x"59D255DD",
x"58AE55C0",
x"57E555CA",
x"57965601",
x"57CF566B",
x"58975708",
x"59DE57CD",
x"5B8A58B2",
x"5D7859A4",
x"5F7C5A92",
x"616F5B69",
x"632E5C1A",
x"64A35C9A",
x"65BB5CE4",
x"667A5CFA",
x"66E95CE3",
x"67165CAC",
x"67195C63",
x"67065C1B",
x"66EF5BE0",
x"66E45BBF",
x"66E65BBF",
x"66FC5BE0",
x"671B5C1C",
x"673F5C6E",
x"67605CC8",
x"67785D1E",
x"677F5D66",
x"67795D97",
x"67685DAC",
x"67545DA7",
x"67445D8A",
x"673E5D5D",
x"674B5D2B",
x"676E5CFB",
x"67A55CD7",
x"67EF5CC6",
x"68455CCB",
x"68A15CE6",
x"68FB5D14",
x"694B5D52",
x"698F5D9A",
x"69C25DE6",
x"69E95E2F",
x"6A0A5E73",
x"6A2B5EAB",
x"6A585ED7",
x"6A975EF4",
x"6AF25F00",
x"6B6B5EFA",
x"6C005EE3",
x"6CAD5EBC",
x"6D625E87",
x"6E105E46",
x"6EA55E00",
x"6F0F5DB6",
x"6F3E5D73",
x"6F275D38",
x"6EC75D0A",
x"6E235CED",
x"6D475CE0",
x"6C455CE6",
x"6B355CFD",
x"6A2E5D22",
x"69475D59",
x"688D5D9F",
x"680A5DF7",
x"67C45E62",
x"67B15EDD",
x"67C85F6A",
x"67FA6000",
x"68376098",
x"68706124",
x"689E6198",
x"68BA61E6",
x"68C56203",
x"68C761E6",
x"68CB6190",
x"68DC6107",
x"6907605A",
x"69585F9A",
x"69D25EDD",
x"6A775E38",
x"6B445DBC",
x"6C2D5D77",
x"6D245D6D",
x"6E1D5D9A",
x"6F025DF6",
x"6FC55E6E",
x"70585EF4",
x"70B15F76",
x"70CC5FE3",
x"70AA6033",
x"704C605F",
x"6FBE6066",
x"6F09604B",
x"6E386015",
x"6D595FCB",
x"6C755F74",
x"6B945F15",
x"6ABD5EB1",
x"69F25E49",
x"69345DDD",
x"68855D6A",
x"67E25CEE",
x"674E5C69",
x"66C85BDA",
x"66545B43",
x"65F55AAC",
x"65AD5A1A",
x"65825995",
x"65755929",
x"658658DA",
x"65B158AE",
x"65F058A5",
x"663558BA",
x"667258E6",
x"6693591A",
x"66835945",
x"66335956",
x"6592593F",
x"649758F4",
x"6342586D",
x"619D57AC",
x"5FB856B9",
x"5DB055A2",
x"5BA3547D",
x"59B85360",
x"58125266",
x"56CF51A5",
x"560C5130",
x"55D45115",
x"562C5158",
x"570D51F7",
x"586552E8",
x"5A1C541B",
x"5C135577",
x"5E2B56E3",
x"60455845",
x"62455981",
x"64175A82",
x"65A95B39",
x"66F35B9B",
x"67F55BA9",
x"68AE5B6B",
x"692B5AF3",
x"69775A55",
x"699E59AF",
x"69B2591B",
x"69BE58B2",
x"69CE5885",
x"69E858A1",
x"6A135904",
x"6A4C59A8",
x"6A905A7A",
x"6ADB5B63",
x"6B235C4D",
x"6B635D24",
x"6B9A5DD2",
x"6BC85E52",
x"6BF55E9E",
x"6C265EC1",
x"6C695EC2",
x"6CC95EB3",
x"6D515EA7",
x"6E045EA7",
x"6EE25EBC",
x"6FE25EEA",
x"70F95F31",
x"72135F84",
x"731D5FDD",
x"74006031",
x"74AF6073",
x"752060A1",
x"754E60B8",
x"753F60BC",
x"750260B2",
x"74A760A5",
x"7442609D",
x"73E8609F",
x"73A760B4",
x"738E60DA",
x"73A06110",
x"73D9614E",
x"7437618E",
x"74AB61CB",
x"752E61FC",
x"75B46222",
x"7638623C",
x"76B56250",
x"77306266",
x"77AB6284",
x"782D62B5",
x"78B862FD",
x"79516360",
x"79F363DA",
x"7A966468",
x"7B2B64FA",
x"7BA7658A",
x"7BF46609",
x"7C09666C",
x"7BDB66AD",
x"7B6966C9",
x"7ABB66C4",
x"79DF66A1",
x"78EB666C",
x"77F66630",
x"771A65F3",
x"766965BF",
x"75F36595",
x"75BC6575",
x"75BF6559",
x"75EF653A",
x"7638650D",
x"768764CE",
x"76C46474",
x"76DF6401",
x"76CB637C",
x"768462E9",
x"76116259",
x"757C61D9",
x"74D16179",
x"74216143",
x"737D6141",
x"72F26172",
x"728461CF",
x"723A624F",
x"720E62DD",
x"71FC6368",
x"71F963D9",
x"71FC641E",
x"71FC642A",
x"71EF63F4",
x"71D16380",
x"719E62D6",
x"71586206",
x"71006122",
x"70996045",
x"702A5F81",
x"6FB55EE9",
x"6F445E86",
x"6ED55E59",
x"6E6A5E5C",
x"6E045E80",
x"6D9D5EAF",
x"6D2A5ED5",
x"6CA05ED7",
x"6BF35EA7",
x"6B165E39",
x"69FD5D8B",
x"68A35CA5",
x"67045B92",
x"652D5A69",
x"6328593B",
x"61105821",
x"5F025729",
x"5D1E5663",
x"5B8555D4",
x"5A51557F",
x"59995561",
x"59685574",
x"59C255B3",
x"5A9F5618",
x"5BEE569F",
x"5D995745",
x"5F865805",
x"619D58DD",
x"63C559C9",
x"65EE5AC2",
x"68065BBF",
x"6A075CB8",
x"6BE95DA2",
x"6DAD5E76",
x"6F4F5F2C",
x"70D25FC6",
x"72356043",
x"737A60AD",
x"74A16107",
x"75AA615F",
x"769461BB",
x"7763621F",
x"781A6290",
x"78BC6307",
x"794C637F",
x"79CF63ED",
x"7A45644B",
x"7AB1648D",
x"7B1364B1",
x"7B6A64B4",
x"7BB9649B",
x"7C00646D",
x"7C3C6434",
x"7C6F63F9",
x"7C9963C5",
x"7CBA639E",
x"7CCF6386",
x"7CD6637D",
x"7CCE6381",
x"7CB16390",
x"7C7D63A3",
x"7C2F63B9",
x"7BCC63D6",
x"7B5963FA",
x"7AE0642B",
x"7A6F646F",
x"7A1664C8",
x"79E2653A",
x"79E265BF",
x"7A1D6656",
x"7A9466F0",
x"7B446781",
x"7C1D67FC",
x"7D0D6852",
x"7DFF6879",
x"7ED9686D",
x"7F87682D",
x"7FF967C2",
x"80246737",
x"8006669D",
x"7FA76607",
x"7F116587",
x"7E58652D",
x"7D906504",
x"7CCF6514",
x"7C27655C",
x"7BA865D8",
x"7B5E667C",
x"7B48673B",
x"7B686806",
x"7BB168CE",
x"7C176984",
x"7C8B6A1E",
x"7CFC6A94",
x"7D5B6AE2",
x"7D986B09",
x"7DB16B09",
x"7DA16AE8",
x"7D6C6AAB",
x"7D196A59",
x"7CB269F3",
x"7C45697F",
x"7BD868FC",
x"7B76686C",
x"7B2067D1",
x"7AD3672D",
x"7A8E6681",
x"7A4865D8",
x"79F76534",
x"799764A1",
x"79226427",
x"789B63CB",
x"7806638E",
x"776D6374",
x"76DC6374",
x"765F638A",
x"760063A8",
x"75C663C6",
x"75B263D9",
x"75C163DA",
x"75E863C8",
x"761E63A1",
x"7654636A",
x"767C632B",
x"769062EA",
x"768962AD",
x"76686276",
x"7631624B",
x"75EF6228",
x"75A8620E",
x"756961FA",
x"753A61E9",
x"751D61D9",
x"751361CC",
x"751461C2",
x"751461BB",
x"750761B9",
x"74DC61B8",
x"748261B4",
x"73E961A4",
x"73076180",
x"71D9613C",
x"705F60CF",
x"6EA06032",
x"6CAB5F63",
x"6A945E66",
x"68725D41",
x"66615C04",
x"64765ABD",
x"62CC5982",
x"61765864",
x"607F5771",
x"5FEE56B5",
x"5FC25636",
x"5FF555F4",
x"607955ED",
x"613E561B",
x"62335674",
x"634456F0",
x"64635785",
x"6586582F",
x"66A358E6",
x"67B559A6",
x"68BD5A6E",
x"69BA5B3D",
x"6AB15C12",
x"6BA35CEA",
x"6C915DC5",
x"6D7D5E9F",
x"6E665F74",
x"6F48603F",
x"702460F9",
x"70F9619D",
x"71C76227",
x"728E6294",
x"735362E4",
x"741A631A",
x"74E56339",
x"75B5634E",
x"768D635C",
x"7769636F",
x"7845638B",
x"791863B5",
x"79DB63EA",
x"7A84642A",
x"7B0A6468",
x"7B66649D",
x"7B9464BF",
x"7B9364C6",
x"7B6564AF",
x"7B16647D",
x"7AB16435",
x"7A4963E5",
x"79F0639B",
x"79BC636C",
x"79BF6365",
x"7A076393",
x"7A9E63FA",
x"7B83649D",
x"7CAA656F",
x"7E036665",
x"7F72676B",
x"80D8686F",
x"8210695E",
x"83006A2B",
x"83916ACF",
x"83B76B45",
x"83766B92",
x"82DE6BBD",
x"820B6BCF",
x"81276BD7",
x"80556BDB",
x"7FBF6BE5",
x"7F836BF8",
x"7FB16C16",
x"804C6C3E",
x"81496C69",
x"828D6C96",
x"83F26CBB",
x"854F6CD4",
x"867D6CDC",
x"875B6CD1",
x"87D26CB1",
x"87D86C7C",
x"876F6C34",
x"86AA6BE1",
x"859E6B87",
x"84696B31",
x"832A6AE6",
x"81FA6AAE",
x"80EF6A8F",
x"80146A8A",
x"7F6C6A9D",
x"7EF36AC1",
x"7E9B6AEB",
x"7E586B0D",
x"7E166B19",
x"7DC66B00",
x"7D606AB8",
x"7CDE6A3E",
x"7C426990",
x"7B9668B7",
x"7AE867BC",
x"7A4966B4",
x"79CF65AD",
x"798764BA",
x"797D63E6",
x"79B5633F",
x"7A2862C9",
x"7ACB6286",
x"7B866270",
x"7C426281",
x"7CE562AF",
x"7D5662EF",
x"7D866334",
x"7D6A6374",
x"7D0663A8",
x"7C6263C9",
x"7B9063D5",
x"7AA463C8",
x"79B563A7",
x"78D56376",
x"780E6339",
x"776262FA",
x"76CC62BB",
x"763B6280",
x"759B6246",
x"74D66209",
x"73D361BE",
x"7286615A",
x"70E260CF",
x"6EE96010",
x"6CA85F14",
x"6A375DD9",
x"67B05C66",
x"65355AC6",
x"62EC5911",
x"60F55764",
x"5F6E55DE",
x"5E69549C",
x"5DF353BC",
x"5E0D534D",
x"5EB3535A",
x"5FD153E0",
x"615654D1",
x"63285618",
x"652E5797",
x"674E5930",
x"69755AC9",
x"6B905C48",
x"6D965D9E",
x"6F7F5EC2",
x"714B5FB7",
x"72FD6081",
x"749E6131",
x"763461D2",
x"77C56272",
x"7958631D",
x"7AEC63D6",
x"7C8164A0",
x"7E116575",
x"7F94664F",
x"80FE6725",
x"824867F2",
x"836968AB",
x"845C6952",
x"851D69E5",
x"85B16A68",
x"861E6ADE",
x"866A6B4E",
x"86A26BBA",
x"86CD6C20",
x"86F96C82",
x"872A6CD7",
x"87656D1A",
x"87AB6D44",
x"88006D4F",
x"885D6D3A",
x"88C26D02",
x"89296CAB",
x"89906C41",
x"89F26BCE",
x"8A4C6B5C",
x"8A9D6AFD",
x"8AE26ABB",
x"8B1A6AA0",
x"8B466AB2",
x"8B676AF7",
x"8B806B69",
x"8B976C06",
x"8BAE6CC2",
x"8BCF6D93",
x"8BFE6E6E",
x"8C436F44",
x"8CA2700A",
x"8D1D70B7",
x"8DAE7145",
x"8E5071B1",
x"8EFD71FB",
x"8FA77226",
x"90427236",
x"90C57234",
x"91277227",
x"91667217",
x"9183720C",
x"91847209",
x"91717212",
x"91567223",
x"913B723D",
x"91277257",
x"911B726A",
x"9117726C",
x"9114725A",
x"91077229",
x"90E771D7",
x"90AB7165",
x"904D70D8",
x"8FCD7037",
x"8F2F6F92",
x"8E7D6EF6",
x"8DC56E76",
x"8D146E1E",
x"8C776DFA",
x"8BF96E0F",
x"8B986E59",
x"8B586ED1",
x"8B2E6F65",
x"8B107003",
x"8AF07093",
x"8AC87105",
x"8A8E714A",
x"8A45715B",
x"89F3713D",
x"89A570F9",
x"896C70A4",
x"895A7054",
x"8980701D",
x"89E67012",
x"8A8E703B",
x"8B737099",
x"8C817123",
x"8DA071C3",
x"8EAE725F",
x"8F8D72DC",
x"90227323",
x"905A731F",
x"902F72C7",
x"8FA57223",
x"8ED27143",
x"8DD3703D",
x"8CCD6F34",
x"8BE56E45",
x"8B366D8C",
x"8AD56D17",
x"8ABE6CEE",
x"8ADD6D02",
x"8B0D6D3E",
x"8B186D7D",
x"8AC56D9A",
x"89D56D6B",
x"88176CCD",
x"856C6BA7",
x"81CB69F0",
x"7D4467B0",
x"780664FA",
x"725161F3",
x"6C765EC6",
x"66CC5BA5",
x"61A758C0",
x"5D4E5640",
x"59F35446",
x"57B352E7",
x"568C522C",
x"566B520F",
x"57265282",
x"5886536E",
x"5A5454B6",
x"5C54563D",
x"5E5757E3",
x"603A598E",
x"61EB5B24",
x"63635C92",
x"64AD5DCD",
x"65D95ED0",
x"67025F98",
x"683E602B",
x"69A36091",
x"6B3860D9",
x"6D006110",
x"6EF3613F",
x"70FD6174",
x"730461B5",
x"74F06203",
x"76A4625C",
x"781062BB",
x"79256314",
x"79E56360",
x"7A556397",
x"7A8663B2",
x"7A8D63B1",
x"7A836397",
x"7A7D636F",
x"7A8D6342",
x"7AC1631F",
x"7B1A6313",
x"7B966325",
x"7C2A6359",
x"7CC963AF",
x"7D62641D",
x"7DE8649A",
x"7E4C6517",
x"7E8B6584",
x"7EA465DB",
x"7E9B6610",
x"7E7D6625",
x"7E596620",
x"7E3F660D",
x"7E4465FA",
x"7E7365FA",
x"7EDB661B",
x"7F7D666A",
x"805B66EF",
x"816A67A7",
x"829D688A",
x"83E3698D",
x"85276A9A",
x"86526BA0",
x"87566C87",
x"88216D3F",
x"88AA6DBD",
x"88ED6DF6",
x"88EC6DEE",
x"88AA6DA4",
x"88326D27",
x"87906C82",
x"86CD6BC5",
x"85FA6B02",
x"85216A47",
x"844F69A1",
x"838E691D",
x"82E968C2",
x"82686893",
x"82106891",
x"81E568B8",
x"81E56900",
x"8209695E",
x"824569C2",
x"828E6A21",
x"82D36A6B",
x"83036A94",
x"83106A96",
x"82EF6A6B",
x"829D6A19",
x"821769A4",
x"81666919",
x"80966881",
x"7FAF67E9",
x"7EC26758",
x"7DD966D2",
x"7CFC6658",
x"7C2B65E5",
x"7B696572",
x"7AAF64F9",
x"79FA6472",
x"794763DD",
x"7894633C",
x"77E86298",
x"774961FE",
x"76C9617D",
x"76766125",
x"765C6101",
x"7687611B",
x"76FD6174",
x"77B86206",
x"78AB62C4",
x"79C1639D",
x"7ADE647F",
x"7BE66558",
x"7CBE6618",
x"7D4F66B5",
x"7D8E672B",
x"7D7A677A",
x"7D1767A8",
x"7C7767BB",
x"7BAE67BC",
x"7ACC67AE",
x"79E36791",
x"78F96762",
x"78096713",
x"77046699",
x"75D965E2",
x"746C64DF",
x"72A76389",
x"707961D8",
x"6DDF5FD6",
x"6AE35D92",
x"679D5B24",
x"643458AE",
x"60D65653",
x"5DB55436",
x"5AFF527A",
x"58D75133",
x"57575071",
x"56855035",
x"565D5072",
x"56C85116",
x"57AA5207",
x"58DE5323",
x"5A445450",
x"5BBD5573",
x"5D2E5675",
x"5E89574F",
x"5FC157FB",
x"60D8587B",
x"61CB58DA",
x"62A15921",
x"635F595C",
x"640A5995",
x"64AA59D7",
x"65425A26",
x"65D95A85",
x"66725AF1",
x"67115B67",
x"67B85BE3",
x"68695C5C",
x"69235CCC",
x"69DE5D2C",
x"6A975D78",
x"6B455DAC",
x"6BDE5DC8",
x"6C5C5DCD",
x"6CB85DC1",
x"6CF05DA9",
x"6D095D91",
x"6D045D7E",
x"6CEB5D7A",
x"6CC85D8A",
x"6CA45DB1",
x"6C875DED",
x"6C795E39",
x"6C795E90",
x"6C8A5EE7",
x"6CAB5F38",
x"6CDB5F7C",
x"6D175FAF",
x"6D5E5FD3",
x"6DAF5FEC",
x"6E0D6000",
x"6E78601A",
x"6EED6041",
x"6F72607E",
x"6FFF60D8",
x"7091614C",
x"712661D8",
x"71B56273",
x"723B6314",
x"72B263AB",
x"731A642E",
x"73726491",
x"73BA64CB",
x"73F664D9",
x"742B64BC",
x"745F647A",
x"7493641D",
x"74CB63AE",
x"7509633C",
x"755162D5",
x"75A06283",
x"75F7624E",
x"76556239",
x"76BA6246",
x"77216270",
x"778762B1",
x"77EC62FE",
x"78466352",
x"789663A3",
x"78D263EC",
x"78FC642B",
x"790E6460",
x"790D6490",
x"78F764BC",
x"78D664EA",
x"78AE651D",
x"788A6553",
x"7870658D",
x"786665C4",
x"787265F0",
x"7894660D",
x"78C86613",
x"790A65FA",
x"795165C5",
x"79966573",
x"79CF650A",
x"79F66491",
x"7A0A6413",
x"7A0C6398",
x"79FD632B",
x"79E562D2",
x"79CB6293",
x"79B7626D",
x"79AA6263",
x"79A8626F",
x"79AB628B",
x"79AD62B4",
x"79A162E0",
x"797F630B",
x"7938632E",
x"78CB6345",
x"78346349",
x"77796339",
x"76A46313",
x"75C262CF",
x"74E06270",
x"740A61F0",
x"7342614E",
x"72836088",
x"71BF5F9E",
x"70E65E91",
x"6FDF5D64",
x"6E975C1C",
x"6D035AC2",
x"6B24595F",
x"690D5801",
x"66DF56B9",
x"64CD559C",
x"630F54BC",
x"61E2542D",
x"617F5404",
x"620A544D",
x"639A5516",
x"662A5664",
x"699A5832",
x"6DBB5A73",
x"72495D15",
x"76FD5FFC",
x"7B936304",
x"7FCF660B",
x"838768EF",
x"86AA6B8F",
x"89376DD2",
x"8B446FAD",
x"8CF3711D",
x"8E70722D",
x"8FE772F1",
x"917E7383",
x"93507403",
x"956E748D",
x"97D6753B",
x"9A7B761C",
x"9D487737",
x"A0197888",
x"A2D27A03",
x"A5527B99",
x"A77B7D30",
x"A9407EB6",
x"AA958016",
x"AB7A8146",
x"ABFA823C",
x"AC2682F6",
x"AC178378",
x"ABE683CC",
x"ABAC83FA",
x"AB87840F",
x"AB878415",
x"ABBD8418",
x"AC30841F",
x"ACE48432",
x"ADCF8454",
x"AEEA848B",
x"B02884D4",
x"B1748531",
x"B2C3859B",
x"B404860F",
x"B52B868B",
x"B6328705",
x"B715877B",
x"B7D487E9",
x"B872884F",
x"B8FB88AC",
x"B9758907",
x"B9F08962",
x"BA7589C3",
x"BB158A2F",
x"BBD68AA8",
x"BCBF8B2E",
x"BDD38BBE",
x"BF0C8C50",
x"C0608CE0",
x"C1B98D60",
x"C2FF8DC5",
x"C4198E06",
x"C4EA8E18",
x"C5558DF7",
x"C54E8DA1",
x"C4C98D15",
x"C3C98C5C",
x"C2608B7B",
x"C0A38A80",
x"BEB98977",
x"BCC38871",
x"BAE7877B",
x"B94386A2",
x"B7ED85EE",
x"B6EB8564",
x"B63F8502",
x"B5D784C6",
x"B5A284A5",
x"B5848492",
x"B5678485",
x"B535846E",
x"B4E18447",
x"B4678408",
x"B3C983B2",
x"B30C8346",
x"B24082CA",
x"B16D8247",
x"B09C81C3",
x"AFD08146",
x"AF0780D3",
x"AE38806A",
x"AD578008",
x"AC577FA9",
x"AB287F45",
x"A9C37ED4",
x"A8257E51",
x"A6537DBA",
x"A45D7D11",
x"A2567C59",
x"A0597B99",
x"9E817ADD",
x"9CE77A2C",
x"9B9F7993",
x"9AB67915",
x"9A2B78B7",
x"99F17875",
x"99F4784D",
x"9A187833",
x"9A3F781F",
x"9A4A7809",
x"9A2877EA",
x"99CF77BE",
x"9940778B",
x"98937751",
x"97DC771F",
x"973C76FC",
x"96D276F1",
x"96AC7702",
x"96D0772D",
x"972B7767",
x"9798779F",
x"97E277BA",
x"97C6779D",
x"9703772C",
x"9563764B",
x"92BE74EF",
x"8F0E7312",
x"8A6970BE",
x"85046E0D",
x"7F326B21",
x"7958682A",
x"73DE6556",
x"6F2B62D6",
x"6B9460D0",
x"69515F63",
x"68795E9B",
x"69075E78",
x"6AD55EED",
x"6DA45FDF",
x"712B612B",
x"751962AF",
x"7924644B",
x"7D0B65DE",
x"80A1674F",
x"83C66893",
x"866F69A1",
x"889E6A79",
x"8A626B21",
x"8BCB6BA3",
x"8CF06C0C",
x"8DE96C6B",
x"8EC86CCB",
x"8F9D6D3D",
x"90736DC8",
x"91526E76",
x"923B6F48",
x"932F703D",
x"942C714E",
x"95287270",
x"961C7395",
x"96FE74A9",
x"97C5759C",
x"9864765B",
x"98D676DE",
x"9914771B",
x"991D7710",
x"98F076C4",
x"98957641",
x"98147595",
x"977674CA",
x"96C573EE",
x"9611730D",
x"9564722F",
x"94C97152",
x"9448707F",
x"93E76FB3",
x"93AB6EF2",
x"93926E3E",
x"939C6D9E",
x"93C86D1D",
x"94116CC2",
x"94776C99",
x"94F96CA6",
x"959A6CEF",
x"965A6D73",
x"97406E2B",
x"984F6F0D",
x"9984700A",
x"9ADC7112",
x"9C487212",
x"9DB372FB",
x"9F0873C0",
x"A028745B",
x"A0F474C6",
x"A1577501",
x"A1437512",
x"A0B47501",
x"9FB574D7",
x"9E64749F",
x"9CE67467",
x"9B677439",
x"9A17741D",
x"991A741A",
x"988E7431",
x"98837464",
x"98F174A9",
x"99C974FB",
x"9AEA754E",
x"9C2B7599",
x"9D6375D2",
x"9E6C75F4",
x"9F2775FB",
x"9F8075E8",
x"9F6E75C1",
x"9EF4758C",
x"9E1C754E",
x"9CF6750D",
x"9B9274CD",
x"9A05748B",
x"98627441",
x"96B173EB",
x"9501737E",
x"935D72F4",
x"91CC724A",
x"90567180",
x"8F04709D",
x"8DDB6FAB",
x"8CDC6EB8",
x"8C0D6DD4",
x"8B6A6D0D",
x"8AED6C6F",
x"8A8E6BFF",
x"8A416BBE",
x"89F96BA3",
x"89A86BA3",
x"89456BAB",
x"88C86BAD",
x"882B6B94",
x"87726B58",
x"869D6AF0",
x"85B26A5B",
x"84BB699E",
x"83BE68C7",
x"82BF67DF",
x"81C366F9",
x"80CB6620",
x"7FD3655E",
x"7ED564B8",
x"7DC9642D",
x"7CA763B5",
x"7B626346",
x"79F062D3",
x"7849624E",
x"766661AD",
x"744560E4",
x"71E85FF7",
x"6F565EE4",
x"6CA05DB5",
x"69D85C74",
x"67175B33",
x"647D5A02",
x"622758F0",
x"6034580B",
x"5EBF575E",
x"5DDC56F3",
x"5D9956CD",
x"5DF356EE",
x"5EE45751",
x"605A57F0",
x"623758C0",
x"645E59B3",
x"66AA5ABC",
x"68FB5BC9",
x"6B325CCD",
x"6D3D5DBD",
x"6F0C5E91",
x"709D5F45",
x"71F35FDD",
x"731A605F",
x"742460D6",
x"75236150",
x"762461D9",
x"7735627A",
x"785D6335",
x"799A640B",
x"7AE364F3",
x"7C2A65E0",
x"7D6066C1",
x"7E736787",
x"7F556821",
x"7FFF6889",
x"806A68B7",
x"80A168B2",
x"80AE6884",
x"80A1683B",
x"808D67E9",
x"808167A0",
x"808A676C",
x"80AE675B",
x"80EC676D",
x"813967A5",
x"818D67FC",
x"81D66866",
x"820968DC",
x"82206952",
x"821569BF",
x"81F36A1E",
x"81C26A6B",
x"81936AA4",
x"81746ACB",
x"81746AE1",
x"819B6AEB",
x"81E96AEB",
x"82596AE5",
x"82DE6ADE",
x"83686AD9",
x"83E26AD7",
x"843F6AD9",
x"84746AE1",
x"84796AEB",
x"844F6AF2",
x"84006AF3",
x"83956AE6",
x"831E6AC7",
x"82AA6A8D",
x"82426A38",
x"81F069C8",
x"81B7693F",
x"819668A8",
x"8187680D",
x"81846777",
x"818466F6",
x"81846691",
x"817D6652",
x"8170663C",
x"815D664E",
x"814C6683",
x"814266D6",
x"8146673E",
x"815D67B4",
x"818B6830",
x"81D068AB",
x"822B6921",
x"8293698E",
x"830169EF",
x"836A6A41",
x"83C66A82",
x"840A6AAE",
x"842C6AC7",
x"842B6ACB",
x"84046ABE",
x"83B96AA6",
x"83506A87",
x"82CF6A6C",
x"82416A5C",
x"81AD6A61",
x"811D6A7C",
x"80986AB0",
x"80286AF7",
x"7FD26B49",
x"7F976B9A",
x"7F7C6BDB",
x"7F7F6BFF",
x"7F9E6BFA",
x"7FD66BCA",
x"80216B6B",
x"80776AE3",
x"80CE6A3D",
x"811A6987",
x"815368CF",
x"816D6824",
x"81636790",
x"812E671A",
x"80CF66C1",
x"80496684",
x"7FA26658",
x"7EE26634",
x"7E116609",
x"7D3565C9",
x"7C52656C",
x"7B6264E6",
x"7A5F6431",
x"793E6349",
x"77F26235",
x"766F60F9",
x"74B45FA1",
x"72C15E3D",
x"70A85CE6",
x"6E8A5BB3",
x"6C8E5ABF",
x"6AE95A25",
x"69D159FE",
x"69765A5A",
x"6A035B46",
x"6B8E5CBD",
x"6E175EB5",
x"71876113",
x"75B463B4",
x"7A5D6670",
x"7F3C691D",
x"84066B94",
x"887A6DB7",
x"8C676F70",
x"8FB170C0",
x"925571AB",
x"9466724A",
x"960A72BB",
x"97767320",
x"98E0739C",
x"9A79744A",
x"9C66753D",
x"9EB87679",
x"A16E77FB",
x"A47179AD",
x"A79B7B79",
x"AAB67D3D",
x"AD8F7EDB",
x"AFF78035",
x"B1C08139",
x"B2D681DA",
x"B32F8216",
x"B2D781F2",
x"B1EB8181",
x"B09280D7",
x"AEFB800A",
x"AD537F33",
x"ABC97E6B",
x"AA7B7DBD",
x"A9847D3A",
x"A8EE7CE5",
x"A8BF7CC1",
x"A8F47CCA",
x"A9887CFE",
x"AA767D57",
x"ABBD7DD3",
x"AD607E72",
x"AF647F36",
x"B1CD8025",
x"B49E8143",
x"B7D08292",
x"BB518412",
x"BF0485BF",
x"C2BF878B",
x"C64D8964",
x"C9798B35",
x"CC108CE6",
x"CDEA8E5D",
x"CEEF8F8A",
x"CF239063",
x"CE9D90E6",
x"CD8E911D",
x"CC33911D",
x"CAD390FE",
x"C9B490E2",
x"C90E90E0",
x"C9079111",
x"C9A99180",
x"CAE5922D",
x"CC96930D",
x"CE849409",
x"D06D9503",
x"D21295DC",
x"D3419679",
x"D3D896C4",
x"D3CA96B4",
x"D322964E",
x"D20195A0",
x"D09394C5",
x"CF0C93DC",
x"CD9F9304",
x"CC75925B",
x"CBAA91F4",
x"CB4D91D9",
x"CB559207",
x"CBB39272",
x"CC499304",
x"CCF193A4",
x"CD8C9437",
x"CDFB94A5",
x"CE2694DF",
x"CE0494DB",
x"CD929499",
x"CCDA9423",
x"CBEE9386",
x"CAE792D6",
x"C9E3922A",
x"C8FF9193",
x"C85B9122",
x"C80C90E2",
x"C82390D6",
x"C8A790FE",
x"C9959152",
x"CADB91C4",
x"CC5B9244",
x"CDF292C1",
x"CF719328",
x"D0A79368",
x"D1679374",
x"D1899342",
x"D0F192CC",
x"CF929210",
x"CD719111",
x"CAA58FD6",
x"C7518E6A",
x"C3A68CD8",
x"BFD48B2A",
x"BC09896C",
x"B86A87A4",
x"B50785D7",
x"B1E08405",
x"AEDC8225",
x"ABD2802B",
x"A8877E07",
x"A4BF7BA3",
x"A04278F1",
x"9AE675E1",
x"949A726C",
x"8D696E99",
x"857F6A75",
x"7D256620",
x"74BE61C3",
x"6CB85D90",
x"658359BC",
x"5F80567B",
x"5AFC53FA",
x"58245257",
x"570051A0",
x"577651D1",
x"594E52D4",
x"5C3D5487",
x"5FE656B8",
x"63F85935",
x"68235BD0",
x"6C2A5E5D",
x"6FE660BC",
x"734562DC",
x"764664B4",
x"78F76645",
x"7B69679A",
x"7DAF68BB",
x"7FDC69B4",
x"81F76A8D",
x"84076B4B",
x"86046BEC",
x"87E96C6F",
x"89A96CCE",
x"8B3C6D09",
x"8C976D1E",
x"8DB46D12",
x"8E8D6CEC",
x"8F216CB8",
x"8F726C80",
x"8F836C51",
x"8F5C6C33",
x"8F066C2B",
x"8E906C3D",
x"8E0A6C65",
x"8D876C9D",
x"8D1A6CE1",
x"8CD36D26",
x"8CC26D69",
x"8CE96DA7",
x"8D4B6DE1",
x"8DDB6E16",
x"8E8A6E4D",
x"8F436E89",
x"8FEE6ED1",
x"90746F24",
x"90C66F85",
x"90D96FEF",
x"90AC705E",
x"904670C7",
x"8FB77124",
x"8F0D716B",
x"8E5C7193",
x"8DB67199",
x"8D287178",
x"8CB87131",
x"8C6770C7",
x"8C357041",
x"8C1E6FA9",
x"8C1E6F06",
x"8C316E65",
x"8C596DD2",
x"8C976D58",
x"8CF06CFD",
x"8D696CCD",
x"8E066CC8",
x"8EC96CF3",
x"8FB16D4F",
x"90B96DD8",
x"91DD6E89",
x"93116F5B",
x"944D7047",
x"95877141",
x"96B57243",
x"97CC7341",
x"98C87430",
x"999E7506",
x"9A4975B9",
x"9AC27641",
x"9B047695",
x"9B0E76B0",
x"9AE07690",
x"9A81763C",
x"99FB75B6",
x"9962750D",
x"98C57454",
x"983F739F",
x"97E77305",
x"97D0729C",
x"98087274",
x"98937297",
x"996C730B",
x"9A8473C7",
x"9BC574BB",
x"9D0E75D1",
x"9E4576EE",
x"9F4677F4",
x"9FFE78C7",
x"A05A7958",
x"A057799C",
x"9FFD7993",
x"9F5C794E",
x"9E9178E4",
x"9DBC7872",
x"9CFD7818",
x"9C7377F4",
x"9C327819",
x"9C497896",
x"9CB87967",
x"9D767A7B",
x"9E6D7BBA",
x"9F877D06",
x"A0A57E3A",
x"A1AB7F36",
x"A27E7FE3",
x"A30B8032",
x"A340801E",
x"A3147FA8",
x"A27B7EDE",
x"A1717DCA",
x"9FEC7C77",
x"9DE37AEE",
x"9B4F7930",
x"9828773D",
x"946F750C",
x"9028729D",
x"8B6A6FEE",
x"86526D0A",
x"81106A04",
x"7BDB66FF",
x"76F2641E",
x"72976190",
x"6F035F7E",
x"6C625E0D",
x"6ACF5D53",
x"6A4F5D53",
x"6AD75E04",
x"6C445F48",
x"6E6960F6",
x"711362DD",
x"741064D0",
x"773266A5",
x"7A586841",
x"7D6F6993",
x"806C6A9D",
x"83536B6B",
x"862A6C14",
x"88FA6CB3",
x"8BC96D61",
x"8E946E30",
x"91506F2B",
x"93EF7054",
x"965571A0",
x"986C72FE",
x"9A1C7455",
x"9B57758D",
x"9C17768D",
x"9C5D7743",
x"9C39779F",
x"9BC0779B",
x"9B0D7739",
x"9A3B767F",
x"9960757E",
x"988D7448",
x"97CA72F6",
x"9718719F",
x"966E705C",
x"95C16F43",
x"95016E63",
x"94286DCD",
x"932E6D85",
x"92176D89",
x"90EE6DD4",
x"8FC56E55",
x"8EB26EFE",
x"8DD06FB9",
x"8D327072",
x"8CEA711A",
x"8D0371A1",
x"8D7A7200",
x"8E487234",
x"8F587241",
x"9095722A",
x"91E771FE",
x"933471C5",
x"9469718F",
x"95777166",
x"96567157",
x"97077162",
x"978B7190",
x"97EA71DB",
x"98287240",
x"984C72B4",
x"9858732F",
x"984A73A3",
x"98257409",
x"97E27458",
x"9784748F",
x"971074AF",
x"969074BD",
x"961174C8",
x"95AB74DB",
x"95737506",
x"957A7554",
x"95D375CB",
x"9684766B",
x"978A772C",
x"98D477FF",
x"9A4C78D3",
x"9BD0798C",
x"9D3C7A18",
x"9E6E7A63",
x"9F497A5E",
x"9FB67A06",
x"9FAC7961",
x"9F2C7878",
x"9E427760",
x"9CFE762A",
x"9B7A74EF",
x"99CF73C1",
x"981172B0",
x"965671C4",
x"94AA7105",
x"9315706F",
x"919B7000",
x"903F6FB3",
x"8F006F7F",
x"8DE06F5E",
x"8CE26F4D",
x"8C0A6F48",
x"8B606F4E",
x"8AEC6F5E",
x"8AB26F78",
x"8AB66F9C",
x"8AF76FC8",
x"8B6D6FFA",
x"8C0D7030",
x"8CC57064",
x"8D867090",
x"8E3970B0",
x"8ED370C1",
x"8F4670BE",
x"8F8870A9",
x"8F9D707F",
x"8F837043",
x"8F416FF9",
x"8EDA6FA6",
x"8E556F48",
x"8DAC6EE2",
x"8CD86E70",
x"8BCB6DEB",
x"8A706D48",
x"88B76C7D",
x"868D6B7F",
x"83E76A45",
x"80C868CC",
x"7D386717",
x"79536532",
x"753E632F",
x"71286128",
x"6D425F38",
x"69C05D7B",
x"66CB5C0D",
x"64845AFD",
x"62FD5A52",
x"62385A0A",
x"622B5A18",
x"62BB5A67",
x"63CA5AE0",
x"65335B67",
x"66D45BEA",
x"68905C59",
x"6A525CAC",
x"6C0D5CEA",
x"6DBF5D1E",
x"6F6B5D57",
x"71165DAB",
x"72CC5E28",
x"74945EE0",
x"76725FD6",
x"78606108",
x"7A5D626D",
x"7C5E63F7",
x"7E536590",
x"80356724",
x"81FC68A3",
x"83A269FC",
x"852C6B2A",
x"86A26C2A",
x"88106D00",
x"89816DB5",
x"8B036E55",
x"8C9B6EE9",
x"8E4F6F7C",
x"90147016",
x"91E270B9",
x"939F7165",
x"953B7217",
x"969A72CA",
x"97A57376",
x"98507416",
x"989374A1",
x"986D7513",
x"97F0756B",
x"972F75A6",
x"964875C7",
x"955D75D1",
x"949275CA",
x"940A75B9",
x"93DF75A5",
x"94257593",
x"94E9758F",
x"9627759C",
x"97D375C0",
x"99D575FC",
x"9C107651",
x"9E5C76BC",
x"A0947736",
x"A29577BA",
x"A442783D",
x"A58478B7",
x"A652791F",
x"A6AF7971",
x"A6A979A6",
x"A65779C1",
x"A5D479C4",
x"A53F79B4",
x"A4B57998",
x"A44A7978",
x"A412795B",
x"A40F794A",
x"A4407947",
x"A49C7956",
x"A5157977",
x"A59C79A6",
x"A62379E1",
x"A69E7A23",
x"A7077A65",
x"A75A7AA3",
x"A79B7ADA",
x"A7CD7B09",
x"A7F87B33",
x"A8217B60",
x"A84F7B95",
x"A8857BDE",
x"A8C77C46",
x"A9147CD1",
x"A9677D85",
x"A9BC7E5D",
x"AA087F49",
x"AA43803A",
x"AA5D8116",
x"AA4A81C2",
x"A9FB8221",
x"A966821E",
x"A88181A9",
x"A74F80C3",
x"A5D67F74",
x"A4287DD4",
x"A25D7BFE",
x"A0957A1C",
x"9EF37853",
x"9D9576C3",
x"9C957589",
x"9C0174B3",
x"9BD77441",
x"9C0D7429",
x"9C847452",
x"9D1774A6",
x"9D9B7505",
x"9DE97554",
x"9DE0757E",
x"9D6D7576",
x"9C8A753B",
x"9B3F74D0",
x"99A27440",
x"97CF7396",
x"95E072DE",
x"93ED7221",
x"91FE715E",
x"9010708F",
x"8E116FA9",
x"8BE56E9C",
x"896A6D58",
x"86876BD2",
x"832A6A06",
x"7F5667F7",
x"7B2365B8",
x"76C26363",
x"7275611A",
x"6E8F5F06",
x"6B5E5D4B",
x"692D5C0E",
x"68355B67",
x"68935B64",
x"6A445C06",
x"6D2A5D3F",
x"710D5EF8",
x"75A16117",
x"7A936377",
x"7F8E65F9",
x"844C687D",
x"88956AEC",
x"8C466D33",
x"8F526F47",
x"91C07123",
x"93A872C4",
x"9529742F",
x"9667756B",
x"97887682",
x"98AE777E",
x"99ED786D",
x"9B5A7958",
x"9CFD7A4A",
x"9ED37B49",
x"A0D67C54",
x"A2F77D6A",
x"A5237E7F",
x"A7437F82",
x"A93F8067",
x"AB008118",
x"AC718188",
x"AD8581AD",
x"AE338188",
x"AE7E811F",
x"AE6B8082",
x"AE097FC3",
x"AD6B7EFA",
x"ACA87E39",
x"ABD27D8F",
x"AAF77D05",
x"AA267C9C",
x"A9667C4A",
x"A8B57C06",
x"A8117BC3",
x"A7757B75",
x"A6DC7B16",
x"A6427AA8",
x"A5A57A2F",
x"A50579B9",
x"A4677954",
x"A3CF7910",
x"A33D78F7",
x"A2B57909",
x"A2307947",
x"A1AB79A5",
x"A11C7A11",
x"A07D7A77",
x"9FC37AC4",
x"9EEC7AE8",
x"9DF87ADA",
x"9CF37A96",
x"9BE77A22",
x"9AE9798B",
x"9A0E78E2",
x"996A783D",
x"991277AD",
x"99127744",
x"996D770F",
x"9A217713",
x"9B257750",
x"9C6777C0",
x"9DD5785A",
x"9F597912",
x"A0DF79DB",
x"A2557AAA",
x"A3AB7B77",
x"A4D77C36",
x"A5CF7CE3",
x"A6887D7A",
x"A6FF7DF4",
x"A72E7E50",
x"A70E7E88",
x"A6A27E98",
x"A5EE7E7C",
x"A4FE7E35",
x"A3E37DBF",
x"A2B27D1E",
x"A1877C5B",
x"A0777B7F",
x"9F9B7A9C",
x"9EFD79BE",
x"9EA178F9",
x"9E7E7858",
x"9E8377E5",
x"9E9477A5",
x"9E977793",
x"9E7477AC",
x"9E1E77DE",
x"9D927820",
x"9CDD7861",
x"9C157896",
x"9B5D78BA",
x"9AD778CA",
x"9AA278C8",
x"9AD578BD",
x"9B7178B0",
x"9C6C78AA",
x"9DA878AD",
x"9EFA78BD",
x"A03378D6",
x"A12478EE",
x"A1A578FF",
x"A19F78FF",
x"A10E78E5",
x"9FFB78AF",
x"9E84785A",
x"9CCC77EB",
x"9AF77762",
x"992576C4",
x"97647610",
x"95B37540",
x"94007447",
x"92227317",
x"8FEE719C",
x"8D366FC3",
x"89D56D83",
x"85B56ADB",
x"80DD67D5",
x"7B6F648D",
x"75A4612B",
x"6FCA5DDF",
x"6A3E5ADF",
x"6559585D",
x"616F5684",
x"5EB85570",
x"5D585528",
x"5D4B55A3",
x"5E7856C4",
x"60A75867",
x"63945A57",
x"66F05C6A",
x"6A705E73",
x"6DD56050",
x"70ED61F2",
x"739B634C",
x"75D66465",
x"77A16542",
x"790C65F3",
x"7A2F6684",
x"7B2166FD",
x"7BF76763",
x"7CC467BA",
x"7D8E67FC",
x"7E5D6828",
x"7F2E683C",
x"8000683B",
x"80CB6826",
x"81886804",
x"823167DF",
x"82BC67C1",
x"832467B1",
x"836267B5",
x"836F67CE",
x"834867F9",
x"82E96830",
x"82566869",
x"8196689D",
x"80AF68C1",
x"7FAF68CF",
x"7EA468C5",
x"7D9D68A0",
x"7CA76865",
x"7BCC6819",
x"7B1667C4",
x"7A84676C",
x"7A1A6719",
x"79D266CF",
x"79A76693",
x"79946663",
x"79936641",
x"799D6627",
x"79AF6613",
x"79C96600",
x"79E965EC",
x"7A0E65D6",
x"7A3865BF",
x"7A6865A7",
x"7A9B6591",
x"7AD26581",
x"7B07657A",
x"7B39657A",
x"7B666583",
x"7B896591",
x"7BA165A3",
x"7BB165B4",
x"7BB965C2",
x"7BBF65CC",
x"7BCB65D2",
x"7BE365D8",
x"7C0E65E0",
x"7C5865F5",
x"7CC46616",
x"7D53664C",
x"7E0A669A",
x"7EE066FF",
x"7FD16779",
x"80CF6804",
x"81D06899",
x"82C96931",
x"83AF69C5",
x"847A6A4E",
x"85276AC5",
x"85B56B2A",
x"86286B76",
x"86876BAA",
x"86D66BC4",
x"871A6BC5",
x"87566BB0",
x"878A6B84",
x"87AF6B45",
x"87BF6AF5",
x"87B16A9A",
x"877C6A37",
x"871A69D1",
x"868B696D",
x"85D66916",
x"850768CC",
x"842F6899",
x"8365687F",
x"82BC6883",
x"824968A7",
x"821868E6",
x"822E693E",
x"828369A7",
x"83096A16",
x"83AA6A7F",
x"844B6AD4",
x"84D06B07",
x"85226B11",
x"85346AEC",
x"84FB6A96",
x"84816A14",
x"83D26972",
x"830668BE",
x"8235680A",
x"81796765",
x"80E566DE",
x"8080667A",
x"8049663E",
x"80316620",
x"80176610",
x"7FD665F9",
x"7F4265C1",
x"7E2D654C",
x"7C6D6486",
x"79E9635C",
x"769461C8",
x"72775FCC",
x"6DAE5D7A",
x"686D5AEB",
x"62F75843",
x"5D9A55AC",
x"58AA534D",
x"54755150",
x"513E4FD3",
x"4F364EEC",
x"4E714EA5",
x"4EEF4EFA",
x"50944FD8",
x"532D512B",
x"567852CE",
x"5A2A54A2",
x"5DFD5682",
x"61AB5853",
x"650359FE",
x"67DF5B74",
x"6A305CAC",
x"6BF55DA8",
x"6D385E69",
x"6E145EF6",
x"6E9E5F58",
x"6EF35F97",
x"6F255FBC",
x"6F455FCF",
x"6F5E5FD9",
x"6F725FE0",
x"6F835FF0",
x"6F93600D",
x"6FA06042",
x"6FAE6090",
x"6FBE60F9",
x"6FD26179",
x"6FF06204",
x"70196290",
x"704A630A",
x"707F6362",
x"70B46387",
x"70E16373",
x"70FD631F",
x"71036291",
x"70ED61D3",
x"70BC60F6",
x"7075600A",
x"701A5F27",
x"6FB55E59",
x"6F4E5DAF",
x"6EEB5D2F",
x"6E945CDA",
x"6E4E5CAF",
x"6E1A5CA7",
x"6DF85CBD",
x"6DE95CED",
x"6DEE5D32",
x"6E035D8E",
x"6E2A5DFE",
x"6E605E86",
x"6EA35F1E",
x"6EF05FC8",
x"6F416077",
x"6F8F6124",
x"6FCF61BF",
x"6FFA6241",
x"700A629B",
x"6FF962C9",
x"6FC862CB",
x"6F7962A4",
x"6F16625F",
x"6EA76206",
x"6E3A61A9",
x"6DD86155",
x"6D8A6114",
x"6D5860EC",
x"6D3F60E0",
x"6D3F60EC",
x"6D55610B",
x"6D796135",
x"6DA56164",
x"6DD96191",
x"6E1061B8",
x"6E4F61D9",
x"6E9661F3",
x"6EE96209",
x"6F4C621E",
x"6FBF6237",
x"70426250",
x"70D2626F",
x"7169628B",
x"71FF62A5",
x"728E62B7",
x"731162B9",
x"738462AB",
x"73E36287",
x"742E624F",
x"74666206",
x"748A61AE",
x"749B614C",
x"749660EA",
x"747A6090",
x"74446041",
x"73F06004",
x"73805FDD",
x"72F65FCD",
x"72565FD3",
x"71AB5FEE",
x"70FF6018",
x"7062604F",
x"6FE0608E",
x"6F8A60D2",
x"6F656117",
x"6F75615C",
x"6FB761A1",
x"702161E3",
x"70A36224",
x"71286260",
x"719C6298",
x"71E862C8",
x"71FC62ED",
x"71CB6301",
x"71516303",
x"708D62EA",
x"6F8762B2",
x"6E4C6255",
x"6CE861CC",
x"6B656115",
x"69D1602D",
x"68315F10",
x"66895DC5",
x"64D85C50",
x"631C5ABD",
x"6152591C",
x"5F7C577E",
x"5D9C55FA",
x"5BBD54A2",
x"59EC538C",
x"584152C9",
x"56CF525E",
x"55B15251",
x"54FB529B",
x"54BD532F",
x"550253F8",
x"55C854E4",
x"570855D9",
x"58B156C2",
x"5AAB5791",
x"5CDC583A",
x"5F2758C0",
x"616E5925",
x"639A5974",
x"659959BD",
x"675C5A0E",
x"68E15A73",
x"6A245AF3",
x"6B2D5B90",
x"6C035C43",
x"6CB15D01",
x"6D425DB6",
x"6DC15E52",
x"6E355EC2",
x"6EA55EFA",
x"6F105EF6",
x"6F755EB5",
x"6FCE5E45",
x"70145DB5",
x"70415D1A",
x"704B5C8A",
x"70305C18",
x"6FE95BD5",
x"6F7D5BC3",
x"6EF05BE9",
x"6E4E5C39",
x"6DA15CAC",
x"6CFC5D31",
x"6C6B5DB8",
x"6BF95E31",
x"6BAE5E90",
x"6B8C5ECD",
x"6B8E5EE7",
x"6BAD5EDA",
x"6BD95EAE",
x"6C095E67",
x"6C2A5E10",
x"6C355DB2",
x"6C275D59",
x"6C005D11",
x"6BCB5CE6",
x"6B965CE3",
x"6B735D10",
x"6B755D70",
x"6BAB5E03",
x"6C205EC3",
x"6CD65FA5",
x"6DC7609B",
x"6EE36190",
x"70166274",
x"71446335",
x"725263C5",
x"732B6420",
x"73BD6441",
x"73FD642E",
x"73F063F0",
x"739E6393",
x"73186324",
x"727662B2",
x"71CF6246",
x"713861EA",
x"70C461A1",
x"707D6170",
x"706B6153",
x"70876148",
x"70CC614B",
x"71316153",
x"71A6615D",
x"721E6162",
x"72906159",
x"72F06141",
x"733A6113",
x"736960D0",
x"737C607A",
x"73756015",
x"73555FAC",
x"73215F48",
x"72DE5EF3",
x"72905EBB",
x"723F5EA7",
x"71F25EBD",
x"71AA5F01",
x"716C5F6D",
x"713B5FFC",
x"711160A1",
x"70EF614E",
x"70CE61F3",
x"70A66283",
x"707262F0",
x"70306332",
x"6FDC6344",
x"6F7A6323",
x"6F0F62D3",
x"6EA0625F",
x"6E3761D0",
x"6DDB6134",
x"6D916097",
x"6D5C6006",
x"6D385F8A",
x"6D235F2B",
x"6D135EE7",
x"6CFD5EBD",
x"6CD95EA4",
x"6C9E5E91",
x"6C455E77",
x"6BCB5E4C",
x"6B315E04",
x"6A795D9C",
x"69AB5D14",
x"68CE5C70",
x"67EC5BBD",
x"67135B0B",
x"664F5A67",
x"65AD59E6",
x"653A598F",
x"65035971",
x"6514598E",
x"657859E3",
x"66345A69",
x"674B5B17",
x"68BD5BDD",
x"6A835CB2",
x"6C965D8B",
x"6EE85E60",
x"716C5F2E",
x"74145FF7",
x"76D460BF",
x"799B618E",
x"7C62626C",
x"7F206360",
x"81D06474",
x"847065AB",
x"86FE6706",
x"897D6884",
x"8BF06A26",
x"8E5C6BE3",
x"90C36DB7",
x"932E6F9C",
x"959C7188",
x"980F7374",
x"9A857554",
x"9CF7771D",
x"9F5978C6",
x"A19C7A41",
x"A3B27B82",
x"A58A7C81",
x"A7157D36",
x"A84A7DA0",
x"A9287DC1",
x"A9AE7DA3",
x"A9E47D53",
x"A9D77CE1",
x"A9987C60",
x"A9337BE1",
x"A8B67B74",
x"A82B7B26",
x"A7977AFB",
x"A6FA7AF5",
x"A6547B0E",
x"A5A27B3C",
x"A4E17B6F",
x"A4157B9F",
x"A3407BBA",
x"A26B7BB9",
x"A1A27B93",
x"A0F37B4D",
x"A06D7AEB",
x"A0197A78",
x"A0047A03",
x"A02F799F",
x"A0957958",
x"A1307940",
x"A1F3795E",
x"A2CA79B2",
x"A3AB7A39",
x"A4817AE5",
x"A5427BAA",
x"A5EA7C71",
x"A6757D29",
x"A6E97DC4",
x"A74A7E37",
x"A7A57E7E",
x"A8027E9F",
x"A8697E9F",
x"A8DC7E8E",
x"A95B7E77",
x"A9E37E64",
x"AA6A7E5D",
x"AAE67E64",
x"AB4D7E75",
x"AB977E8A",
x"ABBD7E9B",
x"ABBF7E9E",
x"AB9B7E8E",
x"AB567E68",
x"AAF17E30",
x"AA717DEA",
x"A9D47D9B",
x"A91C7D46",
x"A8427CF2",
x"A7437C9C",
x"A61C7C41",
x"A4CC7BDB",
x"A3577B63",
x"A1C67AD0",
x"A0267A20",
x"9E887954",
x"9CFE7871",
x"9B9C7782",
x"9A717696",
x"998575BC",
x"98DD7502",
x"98747476",
x"98437420",
x"983C73FF",
x"984D7412",
x"9869744D",
x"987D74A5",
x"987E7506",
x"98667561",
x"982F75A3",
x"97D975BD",
x"976375A3",
x"96D2754E",
x"962774BB",
x"956973F1",
x"949A72F8",
x"93C071E1",
x"92E070C0",
x"92006FAB",
x"91246EBB",
x"904F6DFF",
x"8F846D83",
x"8EC16D48",
x"8DFC6D4A",
x"8D2A6D73",
x"8C366DAD",
x"8B0B6DD4",
x"89916DCA",
x"87B16D6F",
x"85586CAD",
x"827D6B78",
x"7F2269CC",
x"7B5967BB",
x"773F6559",
x"72FC62C8",
x"6EC1602B",
x"6AC55DAB",
x"673D5B6A",
x"64525987",
x"622A5818",
x"60D65729",
x"605C56BD",
x"60B156CD",
x"61BD574F",
x"63615830",
x"6579595D",
x"67DF5AC2",
x"6A705C4B",
x"6D105DE6",
x"6FA55F86",
x"7220611E",
x"747262A7",
x"76966418",
x"78876570",
x"7A4566AB",
x"7BD167C6",
x"7D2A68C1",
x"7E55699A",
x"7F596A51",
x"803E6AE8",
x"810A6B5F",
x"81CB6BBB",
x"82896C03",
x"834C6C3B",
x"841A6C69",
x"84F46C94",
x"85D66CBD",
x"86B56CE5",
x"87836D09",
x"882F6D20",
x"88AA6D24",
x"88E46D0C",
x"88D36CD2",
x"88746C72",
x"87CC6BEC",
x"86E36B47",
x"85CC6A8D",
x"849A69CB",
x"8360690D",
x"822F685F",
x"811667CC",
x"801D6756",
x"7F4666FF",
x"7E9166C1",
x"7DF9669A",
x"7D7A6683",
x"7D136679",
x"7CC4667C",
x"7C90668B",
x"7C8066AD",
x"7C9B66E0",
x"7CE86728",
x"7D696783",
x"7E1B67E9",
x"7EF76852",
x"7FEA68B0",
x"80E268F7",
x"81C86920",
x"82896923",
x"83136906",
x"835F68CE",
x"836C688C",
x"8341684F",
x"82ED682A",
x"82866827",
x"821D684E",
x"81C2689E",
x"81866911",
x"816A6994",
x"816F6A17",
x"818A6A86",
x"81AF6ACE",
x"81D06AE3",
x"81DF6ABD",
x"81CF6A5C",
x"819B69C8",
x"8142690D",
x"80CB683E",
x"803C676D",
x"7FA466AD",
x"7F0D660E",
x"7E8165A0",
x"7E076568",
x"7DA36568",
x"7D50659B",
x"7D0A65F6",
x"7CC86666",
x"7C7F66D6",
x"7C276730",
x"7BB7675C",
x"7B2B6749",
x"7A8466EF",
x"79C5664C",
x"78F5656A",
x"781D645D",
x"7748633F",
x"767F622E",
x"75CB6146",
x"753160A4",
x"74B46055",
x"7453605F",
x"740D60BC",
x"73DC615D",
x"73BD6227",
x"73A462FC",
x"739163BE",
x"737D6450",
x"736864A1",
x"734C64A3",
x"732B6455",
x"730363BF",
x"72D262EF",
x"729761F7",
x"724B60EE",
x"71EB5FE7",
x"716D5EF1",
x"70CB5E18",
x"6FFC5D64",
x"6EFC5CD5",
x"6DC75C66",
x"6C5F5C14",
x"6AC95BD6",
x"69135BA5",
x"67475B7A",
x"657A5B52",
x"63C15B26",
x"622D5AFA",
x"60D25ACC",
x"5FC15A9E",
x"5F035A70",
x"5E9D5A47",
x"5E8F5A24",
x"5ED55A0B",
x"5F6559FE",
x"60345A01",
x"61335A1A",
x"62545A47",
x"63895A90",
x"64C45AF3",
x"65F95B6D",
x"671D5BFA",
x"68285C92",
x"69115D2B",
x"69D45DB6",
x"6A6D5E2B",
x"6ADB5E80",
x"6B215EAE",
x"6B475EB9",
x"6B535EA5",
x"6B575E7E",
x"6B5F5E55",
x"6B795E36",
x"6BB25E33",
x"6C165E56",
x"6CA75EA4",
x"6D625F1A",
x"6E425FAC",
x"6F3A6050",
x"703860F6",
x"712B618E",
x"7206620D",
x"72BB626C",
x"734462AF",
x"73A062DA",
x"73D362FA",
x"73EC6318",
x"73F46341",
x"73FA6379",
x"740963C4",
x"742B641B",
x"74656479",
x"74B764D3",
x"7521651E",
x"75A06555",
x"76306575",
x"76CB6583",
x"77706589",
x"78206593",
x"78D965AE",
x"799B65E8",
x"7A636645",
x"7B2E66C5",
x"7BF66762",
x"7CB2680D",
x"7D5868B2",
x"7DDF6942",
x"7E3C69A8",
x"7E6C69D6",
x"7E6A69C7",
x"7E3C6979",
x"7DE668F3",
x"7D736841",
x"7CEF6773",
x"7C68669D",
x"7BE865CF",
x"7B7A651B",
x"7B27648D",
x"7AF0642E",
x"7ADB6404",
x"7AE2640D",
x"7B036445",
x"7B3764A7",
x"7B796525",
x"7BBF65B4",
x"7C046641",
x"7C3E66BF",
x"7C68671E",
x"7C796753",
x"7C6D6755",
x"7C3F6724",
x"7BED66C1",
x"7B77663A",
x"7AE0659A",
x"7A2D64F6",
x"79636460",
x"788E63EA",
x"77B8639F",
x"76EB6389",
x"763163A1",
x"759363E2",
x"7517643B",
x"74BE649B",
x"748A64EF",
x"74736523",
x"7473652B",
x"747D6500",
x"748764A4",
x"7483641D",
x"74666379",
x"742862C6",
x"73C56218",
x"733E617E",
x"72946101",
x"71D260A8",
x"71016070",
x"702E6052",
x"6F636042",
x"6EAD6033",
x"6E0D6017",
x"6D895FE2",
x"6D1D5F8B",
x"6CC55F11",
x"6C7C5E78",
x"6C3B5DC8",
x"6BFF5D0D",
x"6BC15C53",
x"6B825BA8",
x"6B3F5B18",
x"6AF75AA6",
x"6AAB5A57",
x"6A565A26",
x"69F65A0B",
x"698359FE",
x"68FB59F6",
x"685E59EA",
x"67B359DC",
x"670459C9",
x"666B59BD",
x"65FF59C3",
x"65E559E9",
x"663B5A3C",
x"67215ACA",
x"68A85B9C",
x"6ADB5CB3",
x"6DAE5E0D",
x"710D5F9D",
x"74D26156",
x"78CF6327",
x"7CD464FC",
x"80AF66C5",
x"843C6873",
x"875C69FD",
x"8A016B5F",
x"8C2A6C96",
x"8DE06DA6",
x"8F356E94",
x"903F6F69",
x"9114702A",
x"91C870E1",
x"9267718F",
x"92FA7239",
x"938372DC",
x"9403737B",
x"9474740C",
x"94D2748D",
x"951A74F8",
x"95457543",
x"9552756B",
x"953E756C",
x"95067548",
x"94A87503",
x"942574A1",
x"937D742F",
x"92B573B7",
x"91D57347",
x"90E472EA",
x"8FF472A9",
x"8F157288",
x"8E567288",
x"8DC972A4",
x"8D7A72D7",
x"8D6D7313",
x"8DA5734E",
x"8E17737C",
x"8EB27396",
x"8F647393",
x"90107374",
x"909D7337",
x"90F172E4",
x"90FA7280",
x"90A97215",
x"8FFC71A7",
x"8EF37140",
x"8D9C70E2",
x"8C0D708D",
x"8A5A7043",
x"88A26FFA",
x"86FD6FB3",
x"85816F62",
x"84416F03",
x"83496E90",
x"829B6E08",
x"82376D66",
x"82136CB1",
x"82236BEC",
x"82566B21",
x"829E6A58",
x"82ED699C",
x"833568F5",
x"836D686D",
x"8390680A",
x"839867CE",
x"838467BB",
x"835867CE",
x"83116803",
x"82B56855",
x"824668C2",
x"81C86941",
x"814169CE",
x"80B76A62",
x"80326AF5",
x"7FBE6B80",
x"7F636BF9",
x"7F2E6C57",
x"7F276C93",
x"7F536CA6",
x"7FB46C8F",
x"80466C4E",
x"81016BED",
x"81DC6B79",
x"82C26AFF",
x"83A26A93",
x"846D6A42",
x"85106A1C",
x"857D6A24",
x"85AF6A5B",
x"85A26ABB",
x"85596B35",
x"84DF6BBD",
x"843C6C3D",
x"83846CAA",
x"82C56CFA",
x"820D6D2A",
x"816C6D3D",
x"80EA6D38",
x"808D6D2A",
x"80556D19",
x"803F6D0F",
x"80466D0D",
x"80626D13",
x"80866D1A",
x"80AA6D19",
x"80C76D04",
x"80D66CD4",
x"80D16C82",
x"80B26C0F",
x"80736B79",
x"80096AC8",
x"7F636A00",
x"7E706921",
x"7D196828",
x"7B3F6711",
x"78CF65CC",
x"75B5644B",
x"71E9627E",
x"6D706060",
x"68655DED",
x"62EF5B32",
x"5D485843",
x"57B75546",
x"528A5266",
x"4E0B4FD0",
x"4A7B4DB0",
x"480C4C2F",
x"46DE4B64",
x"46F24B5A",
x"48364C09",
x"4A7F4D5E",
x"4D934F35",
x"51305162",
x"550D53B9",
x"58EB560B",
x"5C8F5832",
x"5FD25A10",
x"629C5B91",
x"64E15CAF",
x"66A75D6C",
x"68005DD0",
x"69025DF1",
x"69C75DE0",
x"6A665DB6",
x"6AF65D84",
x"6B875D5D",
x"6C215D4C",
x"6CC85D57",
x"6D795D7E",
x"6E305DBB",
x"6EE35E07",
x"6F8C5E56",
x"70215E9F",
x"70A05ED7",
x"71045EFC",
x"714C5F0B",
x"717A5F08",
x"718E5EFD",
x"718D5EEE",
x"71775EE9",
x"71515EF1",
x"71195F0A",
x"70D45F32",
x"707D5F63",
x"70175F97",
x"6FA05FC1",
x"6F135FDA",
x"6E705FDF",
x"6DB85FCF",
x"6CE95FAF",
x"6C0A5F87",
x"6B215F60",
x"6A385F42",
x"695B5F35",
x"68975F38",
x"67FA5F46",
x"67905F55",
x"675E5F58",
x"67605F41",
x"67915F01",
x"67E25E92",
x"683D5DF6",
x"688A5D2E",
x"68B75C4B",
x"68B05B5D",
x"686F5A7B",
x"67F559B9",
x"674E5926",
x"669358CD",
x"65DC58B2",
x"654858D3",
x"64F25929",
x"64EE59AC",
x"65455A4D",
x"65F85B05",
x"66FC5BC9",
x"68405C92",
x"69A85D5D",
x"6B1D5E27",
x"6C875EEC",
x"6DD45FAB",
x"6EF36060",
x"6FDC6107",
x"708D619D",
x"7104621B",
x"71456283",
x"715362D2",
x"7134630A",
x"70EC632E",
x"70866342",
x"700D634B",
x"6F8C634B",
x"6F116345",
x"6EAD6337",
x"6E6F6321",
x"6E5F6300",
x"6E8362D0",
x"6EDE6295",
x"6F656250",
x"700C6207",
x"70C161C1",
x"716F6188",
x"72026168",
x"72686164",
x"72966183",
x"728961C3",
x"7244621D",
x"71CF6284",
x"713A62E9",
x"7099633B",
x"6FFA6369",
x"6F756363",
x"6F136324",
x"6EDC62A8",
x"6ED461F4",
x"6EF56113",
x"6F326014",
x"6F805F0B",
x"6FC85E0A",
x"6FFA5D1F",
x"70035C5A",
x"6FD45BC3",
x"6F625B5C",
x"6EA85B21",
x"6DA45B0A",
x"6C585B0E",
x"6AC85B21",
x"68FB5B31",
x"66F95B32",
x"64C95B1A",
x"62755ADF",
x"60065A7B",
x"5D8859F1",
x"5B0A5943",
x"58A4587B",
x"566B57A5",
x"547956CF",
x"52EE560B",
x"51E25568",
x"516B54F7",
x"519754C0",
x"526C54C9",
x"53DF5512",
x"55DE5595",
x"584A5647",
x"5AFD571C",
x"5DD25801",
x"609D58EB",
x"633B59CC",
x"65935A9E",
x"67945B5D",
x"693B5C0D",
x"6A905CB1",
x"6BA15D53",
x"6C865DFA",
x"6D585EAE",
x"6E2D5F74",
x"6F17604B",
x"70206132",
x"71486222",
x"72896314",
x"73D36400",
x"751764DC",
x"763C65A1",
x"7734664C",
x"77F066DB",
x"7867674B",
x"789B679E",
x"789467D5",
x"785D67F3",
x"780967F7",
x"77A767E6",
x"774567BF",
x"76F06784",
x"76AD673A",
x"767A66DF",
x"7655667A",
x"7635660E",
x"7613659E",
x"75E6652E",
x"75A864C2",
x"755E645A",
x"750763FA",
x"74B163A3",
x"74666358",
x"7437631D",
x"743162F7",
x"746262EF",
x"74D46309",
x"7587634B",
x"767D63B9",
x"77A86456",
x"78FA651B",
x"7A5F65FF",
x"7BBF66F5",
x"7D0067E8",
x"7E0B68C7",
x"7ECE697D",
x"7F3B6A00",
x"7F4F6A44",
x"7F106A47",
x"7E8D6A10",
x"7DDF69AE",
x"7D206932",
x"7C7068B4",
x"7BED6845",
x"7BAE67F7",
x"7BC267D9",
x"7C2D67ED",
x"7CE96832",
x"7DE868A1",
x"7F0D692D",
x"803F69C8",
x"81636A62",
x"825D6AF0",
x"831D6B69",
x"839A6BCA",
x"83D06C12",
x"83CC6C44",
x"83976C65",
x"83446C7C",
x"82DF6C8C",
x"82766C97",
x"82136CA3",
x"81B56CA8",
x"815B6CA8",
x"80FC6C9C",
x"80906C7F",
x"800E6C4E",
x"7F766C04",
x"7EC56BA3",
x"7E016B28",
x"7D356A9A",
x"7C7069FC",
x"7BC26955",
x"7B3768AB",
x"7AD96809",
x"7AAD6775",
x"7AAE66F5",
x"7AD2668D",
x"7B0A6641",
x"7B42660E",
x"7B6365F2",
x"7B5965E8",
x"7B1465E6",
x"7A8A65E5",
x"79B765DB",
x"789D65BF",
x"7746658A",
x"75C46538",
x"742164C2",
x"72726427",
x"70C56368",
x"6F276284",
x"6D9E6183",
x"6C316069",
x"6ADF5F3F",
x"69A75E10",
x"68875CE3",
x"677C5BC9",
x"66875ACD",
x"65AE59FD",
x"64F85966",
x"64725911",
x"642E5905",
x"64415949",
x"64BE59DC",
x"65B85AB8",
x"673D5BDA",
x"69545D38",
x"6BF95EC3",
x"6F236072",
x"72B76235",
x"76966401",
x"7A9865C6",
x"7E93677A",
x"825D6913",
x"85D06A86",
x"88D26BCF",
x"8B526CE9",
x"8D4C6DD7",
x"8EC86E9A",
x"8FD66F3A",
x"90906FC1",
x"910E7039",
x"916A70AD",
x"91B87123",
x"9209719F",
x"92627221",
x"92C972A6",
x"933C7325",
x"93B87393",
x"943C73E8",
x"94C5741D",
x"95537431",
x"95E9742C",
x"96867413",
x"972973F8",
x"97CD73E8",
x"986A73F5",
x"98F67427",
x"99627483",
x"999F7505",
x"99A4759F",
x"996A7640",
x"98F076D0",
x"983E7739",
x"975F776A",
x"96667752",
x"956676F2",
x"9471764D",
x"9398756F",
x"92E6746C",
x"9260735E",
x"9207725B",
x"91D87176",
x"91CA70C0",
x"91D67040",
x"91F16FF9",
x"92136FE5",
x"92346FFA",
x"924F702D",
x"925D7069",
x"925F70A6",
x"924E70D4",
x"922B70EE",
x"91F970EC",
x"91B470D2",
x"916370A1",
x"91067061",
x"909E7016",
x"902E6FCB",
x"8FB56F86",
x"8F346F4E",
x"8EA86F27",
x"8E0E6F13",
x"8D666F0F",
x"8CB16F1C",
x"8BF06F34",
x"8B2E6F52",
x"8A716F73",
x"89C86F92",
x"893C6FA7",
x"88D96FB3",
x"88A76FAE",
x"88A56F9C",
x"88D26F79",
x"89246F47",
x"89906F0A",
x"8A066EC7",
x"8A766E82",
x"8AD26E44",
x"8B106E13",
x"8B2C6DF5",
x"8B246DEE",
x"8AFB6DFF",
x"8AB96E26",
x"8A6A6E5F",
x"8A176EA1",
x"89CB6EE6",
x"89906F23",
x"896D6F4E",
x"89666F64",
x"897C6F61",
x"89A86F45",
x"89E46F14",
x"8A226ED4",
x"8A556E86",
x"8A6A6E33",
x"8A566DDC",
x"8A0E6D85",
x"898E6D2B",
x"88D96CD2",
x"87FE6C79",
x"87126C26",
x"86326BDB",
x"857A6BA6",
x"850A6B8F",
x"84F66BA0",
x"85496BE1",
x"85FE6C52",
x"87046CEC",
x"88346DA1",
x"895C6E57",
x"8A456EEC",
x"8AAF6F41",
x"8A6A6F31",
x"89496EA4",
x"87386D88",
x"84356BDC",
x"805969B0",
x"7BD26721",
x"76E06459",
x"71CF618B",
x"6CF05EEA",
x"68935CA5",
x"64F85AE3",
x"625459BB",
x"60C55939",
x"60545959",
x"60F05A0B",
x"627F5B35",
x"64CD5CB8",
x"67A35E77",
x"6AC76052",
x"6DFC6231",
x"711163FF",
x"73D965A8",
x"76356723",
x"78166860",
x"7972695B",
x"7A4F6A09",
x"7ABE6A69",
x"7AD36A7A",
x"7AAA6A41",
x"7A5C69C8",
x"7A076923",
x"79C16863",
x"799A67A3",
x"799E66FA",
x"79CF6680",
x"7A2A663F",
x"7AA56642",
x"7B316683",
x"7BBF66F6",
x"7C416789",
x"7CA76821",
x"7CEC68AA",
x"7D0A6909",
x"7D016931",
x"7CDA6919",
x"7C9D68BF",
x"7C4F682D",
x"7BFD676D",
x"7BAE6694",
x"7B6665B4",
x"7B2A64DE",
x"7AF9641E",
x"7AD36380",
x"7AB86309",
x"7AA762B8",
x"7AA1628E",
x"7AA46287",
x"7AB5629D",
x"7AD262CC",
x"7AFE6310",
x"7B386365",
x"7B8063C8",
x"7BD36438",
x"7C2F64B1",
x"7C90652F",
x"7CF365AE",
x"7D586627",
x"7DBB6696",
x"7E1E66F2",
x"7E816737",
x"7EE66760",
x"7F4B6772",
x"7FAF676B",
x"80166752",
x"807A6730",
x"80DD6710",
x"813C66FF",
x"819A6706",
x"81F7672D",
x"8259677C",
x"82C567F2",
x"833F688D",
x"83CF6947",
x"84776A17",
x"853B6AF0",
x"86166BC8",
x"87036C93",
x"87F76D48",
x"88E66DDE",
x"89C16E4F",
x"8A776E9A",
x"8AFE6EBA",
x"8B4B6EAE",
x"8B586E79",
x"8B216E1C",
x"8AAB6D9A",
x"89FD6CFA",
x"891F6C45",
x"88216B86",
x"870B6AC8",
x"85EC6A1A",
x"84CF6987",
x"83C1691A",
x"82C968D6",
x"81F268BF",
x"814168CE",
x"80B968F9",
x"80636935",
x"803E6976",
x"804869AE",
x"807D69D5",
x"80D869E6",
x"814869E2",
x"81C369CC",
x"823969B0",
x"82976993",
x"82CE6980",
x"82D0697D",
x"8295698C",
x"821A69A4",
x"815D69C1",
x"806A69D5",
x"7F4B69D1",
x"7E1069A7",
x"7CC8694F",
x"7B8468C1",
x"7A4F67FC",
x"79326703",
x"782D65E0",
x"773A64A0",
x"76506350",
x"75666200",
x"746F60C1",
x"735F5F9E",
x"72355EA4",
x"70F55DDA",
x"6FA85D49",
x"6E635CF1",
x"6D415CD5",
x"6C5B5CF3",
x"6BCF5D46",
x"6BB75DCD",
x"6C275E81",
x"6D285F5D",
x"6EBE605A",
x"70DF6177",
x"737A62AE",
x"767963F9",
x"79BF6555",
x"7D2F66BE",
x"80A8682D",
x"840D699C",
x"87416B02",
x"8A2E6C54",
x"8CC26D89",
x"8EEF6E9A",
x"90AC6F82",
x"91FE7040",
x"92EC70D7",
x"93837151",
x"93D971BB",
x"94067223",
x"94227295",
x"94487319",
x"948673B3",
x"94E6745F",
x"9569750F",
x"960475B4",
x"96A7763A",
x"973B768F",
x"97AB76A6",
x"97E47679",
x"97DA760F",
x"978D7574",
x"970374BE",
x"964D7406",
x"95817365",
x"94B672EE",
x"93FE72A7",
x"93697292",
x"92FB72A0",
x"92B272C0",
x"928472DA",
x"926672D7",
x"924A72A7",
x"92297247",
x"91FE71BA",
x"91CE7114",
x"919D706E",
x"917B6FE5",
x"91716F96",
x"918B6F94",
x"91C96FEB",
x"92287094",
x"929F7182",
x"93217299",
x"939C73B9",
x"940774C1",
x"94567595",
x"948D7622",
x"94AF7662",
x"94CF765E",
x"94FE7625",
x"954D75D2",
x"95D07583",
x"96917554",
x"978E755A",
x"98C075A2",
x"9A15762A",
x"9B7676E8",
x"9CC377C7",
x"9DDF78A7",
x"9EAE796A",
x"9F1979EF",
x"9F117A1F",
x"9E8F79E5",
x"9D9A793D",
x"9C3B782A",
x"9A8776BD",
x"9898750F",
x"968A733E",
x"947D7170",
x"928D6FC3",
x"90CF6E55",
x"8F566D3A",
x"8E2A6C7D",
x"8D466C1D",
x"8CA56C12",
x"8C346C47",
x"8BDA6CA6",
x"8B836D16",
x"8B156D7D",
x"8A846DCB",
x"89C86DF5",
x"88E36DF8",
x"87E36DDC",
x"86E06DAD",
x"85F66D7F",
x"85426D62",
x"84DD6D68",
x"84DA6D9C",
x"853E6E02",
x"86016E93",
x"87116F44",
x"884D7003",
x"899170BB",
x"8AB47155",
x"8B9071C0",
x"8C0B71EE",
x"8C1571DB",
x"8BAC7189",
x"8ADA7103",
x"89B57057",
x"88586F93",
x"86DF6EC8",
x"855F6E02",
x"83E76D44",
x"827A6C8C",
x"81106BCF",
x"7F936B00",
x"7DEC6A0A",
x"7C0068DC",
x"79BA6768",
x"770D65A7",
x"73FC639E",
x"7097615A",
x"6CFD5EF4",
x"695B5C8D",
x"65E15A49",
x"62C5584D",
x"603756B9",
x"5E5C55A8",
x"5D4D5526",
x"5D105533",
x"5DA055C6",
x"5EE456C6",
x"60BB5817",
x"62FB5998",
x"65785B28",
x"680C5CAC",
x"6A905E10",
x"6CEC5F48",
x"6F106052",
x"70F36131",
x"729761F2",
x"740662A1",
x"754C634C",
x"767663FF",
x"779464C1",
x"78B06594",
x"79D16677",
x"7AF66763",
x"7C20684C",
x"7D466928",
x"7E6069E9",
x"7F626A83",
x"80416AEC",
x"80F46B1E",
x"81736B19",
x"81BC6ADF",
x"81CF6A79",
x"81B169F2",
x"816A6959",
x"810668BF",
x"80916837",
x"801A67CE",
x"7FAA6790",
x"7F4B6783",
x"7F0367AA",
x"7ED367FD",
x"7EBE6875",
x"7EBA6903",
x"7EC46999",
x"7ED26A28",
x"7EE36AA3",
x"7EF06B02",
x"7EFD6B3B",
x"7F0B6B52",
x"7F216B45",
x"7F486B19",
x"7F876AD4",
x"7FE26A7A",
x"805B6A11",
x"80ED699E",
x"81906923",
x"823568A1",
x"82CC681E",
x"8345679A",
x"8393671A",
x"83AD66A3",
x"83936638",
x"834C65E0",
x"82E465A1",
x"8273657D",
x"820B6579",
x"81C26594",
x"81AB65D0",
x"81D0662B",
x"823166A3",
x"82C96731",
x"838967D3",
x"84586881",
x"85216934",
x"85C969E5",
x"863E6A87",
x"866F6B13",
x"86536B7F",
x"85ED6BC1",
x"85466BD4",
x"846C6BB7",
x"83736B6B",
x"82706AF7",
x"81776A65",
x"809869C1",
x"7FDF691A",
x"7F4C687C",
x"7EE267F0",
x"7E96677F",
x"7E5D6725",
x"7E3066E2",
x"7E0166AE",
x"7DCF6680",
x"7D986650",
x"7D63661B",
x"7D3865E0",
x"7D2565A3",
x"7D38656A",
x"7D7A653F",
x"7DF0652E",
x"7E97653E",
x"7F656573",
x"804565CE",
x"81226645",
x"81E266CE",
x"826F675C",
x"82B467DE",
x"82AB6846",
x"8252688D",
x"81B268AE",
x"80DF68A8",
x"7FED6884",
x"7EF36849",
x"7E036803",
x"7D2867B8",
x"7C69676D",
x"7BBE6720",
x"7B1866CC",
x"7A686665",
x"799165E0",
x"78866532",
x"77346452",
x"7596633B",
x"73B261F4",
x"71966087",
x"6F595F07",
x"6D1A5D8A",
x"6AFA5C29",
x"69195AFB",
x"67905A15",
x"66735982",
x"65CC594A",
x"659D596A",
x"65D959D7",
x"66735A82",
x"67555B57",
x"68685C43",
x"69965D33",
x"6ACC5E17",
x"6BFD5EE4",
x"6D1D5F95",
x"6E286028",
x"6F1B60A4",
x"6FFC610B",
x"70CB616A",
x"719061C8",
x"724F622B",
x"73116298",
x"73D96311",
x"74AD6397",
x"75936425",
x"768B64B8",
x"77986549",
x"78BC65D5",
x"79F36655",
x"7B3766C6",
x"7C84672A",
x"7DD2677C",
x"7F1A67C1",
x"805667FA",
x"8181682D",
x"829B685E",
x"83A26891",
x"849D68C9",
x"858A690A",
x"86706955",
x"875169A7",
x"88286A02",
x"88F66A5F",
x"89B26ABE",
x"8A556B19",
x"8AD36B6B",
x"8B276BB2",
x"8B4E6BED",
x"8B456C1A",
x"8B136C3D",
x"8AC26C55",
x"8A606C66",
x"89FE6C73",
x"89AE6C82",
x"89816C92",
x"89866CA7",
x"89C56CC1",
x"8A466CE3",
x"8B0A6D0D",
x"8C0D6D41",
x"8D486D7F",
x"8EAC6DC7",
x"902C6E1C",
x"91B26E7A",
x"932A6EE1",
x"947E6F4B",
x"959A6FB3",
x"966E7012",
x"96EE7061",
x"9717709C",
x"96EE70BD",
x"968370C8",
x"95EA70C4",
x"954370B9",
x"94AB70B1",
x"944270BB",
x"941E70E4",
x"944C7130",
x"94CD71A1",
x"95957234",
x"968A72DB",
x"978B7388",
x"98717426",
x"991E74A7",
x"997474FC",
x"9967751D",
x"98F9750C",
x"983674D1",
x"973C7478",
x"96287413",
x"951E73B6",
x"9438736E",
x"93857343",
x"93107337",
x"92C97345",
x"92A17364",
x"927E737E",
x"92457383",
x"91E37365",
x"91497317",
x"90797296",
x"8F7D71E4",
x"8E69710A",
x"8D56701C",
x"8C5D6F2D",
x"8B936E4F",
x"8B046D96",
x"8AAF6D0C",
x"8A8E6CBA",
x"8A8E6C9C",
x"8A9B6CAB",
x"8AA16CD8",
x"8A916D16",
x"8A626D51",
x"8A156D7C",
x"89B56D8F",
x"89506D82",
x"88F66D57",
x"88B76D10",
x"889A6CB5",
x"889D6C4B",
x"88B56BD4",
x"88C86B4C",
x"88B46AB0",
x"885569F0",
x"87806900",
x"861667D3",
x"83FD665F",
x"813164A3",
x"7DBB62A2",
x"79B76072",
x"75555E29",
x"70D25BEE",
x"6C7359E4",
x"68805832",
x"653B56F4",
x"62DB5644",
x"6183562B",
x"614456A5",
x"621957A5",
x"63E65911",
x"66825AC9",
x"69B45CAC",
x"6D415E9A",
x"70ED6076",
x"7483622D",
x"77D963B1",
x"7AD164FD",
x"7D5B6617",
x"7F726704",
x"811D67CF",
x"82686883",
x"83636928",
x"842069C8",
x"84AE6A63",
x"85186AFA",
x"85696B8A",
x"85A56C0D",
x"85CF6C7D",
x"85E96CD8",
x"85F46D19",
x"85F06D3F",
x"85E06D51",
x"85C66D51",
x"85A76D45",
x"85876D3A",
x"856C6D31",
x"855B6D34",
x"85536D42",
x"85586D5C",
x"85656D7C",
x"85746D9C",
x"857F6DB1",
x"857A6DB5",
x"855D6DA3",
x"85206D76",
x"84BC6D30",
x"84316CD4",
x"83806C6B",
x"82B26C00",
x"81D86BA1",
x"80FE6B58",
x"80396B30",
x"7FA06B2D",
x"7F416B55",
x"7F2C6BA7",
x"7F6D6C1E",
x"80096CB4",
x"81006D63",
x"824C6E21",
x"83E56EE6",
x"85BB6FAB",
x"87BB706B",
x"89D3711D",
x"8BEC71C0",
x"8DF07250",
x"8FCC72C7",
x"916F7327",
x"92CA736C",
x"93D67399",
x"949073AD",
x"94F973AD",
x"9518739A",
x"94F67379",
x"94A1734E",
x"9425731A",
x"939172DF",
x"92EF729D",
x"92497252",
x"91A971FC",
x"91187197",
x"909D7123",
x"903C70A1",
x"8FFD7014",
x"8FE06F83",
x"8FEC6EF5",
x"901B6E75",
x"906D6E0A",
x"90D96DBE",
x"91536D97",
x"91CC6D94",
x"92356DB3",
x"927D6DEE",
x"92956E3A",
x"92796E8D",
x"921F6EDE",
x"918E6F20",
x"90CC6F51",
x"8FE66F6C",
x"8EED6F72",
x"8DF06F65",
x"8CFD6F4A",
x"8C206F24",
x"8B596EF6",
x"8AAE6EC3",
x"8A176E8A",
x"898D6E4A",
x"89086E00",
x"88806DAD",
x"87F26D4D",
x"875D6CE3",
x"86C96C76",
x"86426C07",
x"85D96BA3",
x"85A16B51",
x"85B16B1D",
x"86186B0F",
x"86E66B30",
x"881E6B83",
x"89B86C0A",
x"8B9E6CBE",
x"8DB26D94",
x"8FC36E7A",
x"919D6F58",
x"93007013",
x"93B2708A",
x"938170A4",
x"92467048",
x"8FF46F65",
x"8C956DF9",
x"884C6C0C",
x"835969B7",
x"7E0A671B",
x"78BE646A",
x"73D561D6",
x"6FA55F90",
x"6C765DC3",
x"6A755C94",
x"69B25C14",
x"6A245C43",
x"6BA65D15",
x"6E035E6C",
x"70F76021",
x"7444620D",
x"77AB6404",
x"7B0065E9",
x"7E2267A0",
x"81046921",
x"83A86A6C",
x"86186B8D",
x"88666C97",
x"8AA46DA1",
x"8CE36EBF",
x"8F2C7005",
x"91857175",
x"93ED7312",
x"965C74D1",
x"98CA76A0",
x"9B2C786A",
x"9D787A13",
x"9FA57B89",
x"A1A97CB7",
x"A37D7D94",
x"A5187E19",
x"A6757E50",
x"A78F7E41",
x"A8617DFF",
x"A8E97D9B",
x"A9247D2A",
x"A9187CBD",
x"A8CA7C63",
x"A8467C20",
x"A7947BFE",
x"A6C27BF4",
x"A5DC7BFE",
x"A4EC7C12",
x"A3FB7C25",
x"A3127C2D",
x"A2337C20",
x"A1617BFE",
x"A09B7BC1",
x"9FE17B74",
x"9F327B1E",
x"9E8E7ACA",
x"9DF47A89",
x"9D677A68",
x"9CEA7A74",
x"9C827AB3",
x"9C317B25",
x"9BFD7BC6",
x"9BE97C88",
x"9BF37D59",
x"9C1A7E22",
x"9C577ECC",
x"9CA27F40",
x"9CEE7F72",
x"9D2C7F59",
x"9D4F7EF2",
x"9D4B7E47",
x"9D187D6A",
x"9CB67C6F",
x"9C2B7B6F",
x"9B807A82",
x"9AC879B9",
x"9A147923",
x"997978C3",
x"99017898",
x"98B97896",
x"989D78B2",
x"98A578D6",
x"98C378F4",
x"98E278FC",
x"98E978E2",
x"98C878A5",
x"9871783E",
x"97DD77B4",
x"9711770F",
x"961A7655",
x"95077592",
x"93ED74CE",
x"92E47412",
x"91F97362",
x"913872C7",
x"90A47243",
x"903971D7",
x"8FF27188",
x"8FC17157",
x"8F9D7145",
x"8F7D7157",
x"8F5D7189",
x"8F3E71DC",
x"8F24724E",
x"8F1572DA",
x"8F1F7379",
x"8F497425",
x"8F9E74D2",
x"901F7578",
x"90D2760B",
x"91AF7681",
x"92AF76D5",
x"93C87701",
x"94EC7703",
x"960D76DE",
x"971F7696",
x"98177634",
x"98ED75C3",
x"99A1754E",
x"9A3174E2",
x"9AA17488",
x"9AF47446",
x"9B2F741D",
x"9B4F7408",
x"9B4B73F9",
x"9B1773E4",
x"9A9E73B1",
x"99C5734A",
x"9871729C",
x"968B7197",
x"94037037",
x"90D86E7D",
x"8D186C7A",
x"88E66A4B",
x"84766810",
x"800665F5",
x"7BDF6423",
x"784662BF",
x"757A61E8",
x"73AA61AF",
x"72EC6218",
x"73426317",
x"74966497",
x"76BF6675",
x"798A688A",
x"7CBB6AAE",
x"801A6CBD",
x"83776E99",
x"86AF7031",
x"89AB717B",
x"8C637279",
x"8ED97337",
x"911873C7",
x"932E743B",
x"952474AA",
x"97047525",
x"98D475B7",
x"9A947667",
x"9C3D7737",
x"9DD07822",
x"9F46791D",
x"A09C7A1F",
x"A1D37B1B",
x"A2EB7C05",
x"A3EA7CD3",
x"A4D27D7E",
x"A5A57E02",
x"A6677E60",
x"A7197E9B",
x"A7BF7EB7",
x"A8577EC0",
x"A8E67EC1",
x"A9717EC7",
x"AA007EE1",
x"AA987F19",
x"AB457F81",
x"AC0F801C",
x"ACFD80F0",
x"AE0E81F8",
x"AF46832D",
x"B09F847E",
x"B20E85D7",
x"B3888722",
x"B5048846",
x"B6758931",
x"B7D789D6",
x"B9238A31",
x"BA5C8A46",
x"BB818A27",
x"BC9889E4",
x"BDA28997",
x"BEA08959",
x"BF92893C",
x"C06E894D",
x"C129898F",
x"C1B789FE",
x"C20B8A88",
x"C2158B1A",
x"C1CD8B98",
x"C12D8BEF",
x"C03C8C0A",
x"BEFF8BE0",
x"BD8B8B70",
x"BBF78AC2",
x"BA5A89E9",
x"B8D488FE",
x"B77D881B",
x"B669875E",
x"B5A986DE",
x"B54686AF",
x"B53D86D4",
x"B589874F",
x"B61C8811",
x"B6E38907",
x"B7CA8A15",
x"B8C08B21",
x"B9B68C0E",
x"BA9F8CC9",
x"BB778D45",
x"BC398D7D",
x"BCE78D79",
x"BD828D43",
x"BE088CED",
x"BE718C87",
x"BEB28C1E",
x"BEB98BB8",
x"BE708B55",
x"BDBF8AED",
x"BC948A73",
x"BAE189D3",
x"B8A58903",
x"B5EB87F6",
x"B2D086AB",
x"AF7E852B",
x"AC268387",
x"A8FE81D3",
x"A63D802F",
x"A40C7EB5",
x"A2877D77",
x"A1B67C86",
x"A18E7BE8",
x"A1EE7B96",
x"A2A97B85",
x"A3887BA0",
x"A4547BD0",
x"A4DD7BFC",
x"A4FD7C13",
x"A4A17C05",
x"A3C77BC7",
x"A2807B58",
x"A0E77ABC",
x"9F1E79F7",
x"9D497913",
x"9B87781C",
x"99E97719",
x"98707610",
x"97127503",
x"95B373EE",
x"943472CB",
x"92677192",
x"902E703A",
x"8D6C6EBA",
x"8A176D0F",
x"86386B3A",
x"81EC6944",
x"7D65673E",
x"78DF653E",
x"74A16360",
x"70F361C1",
x"6E13607A",
x"6C335FA2",
x"6B6F5F48",
x"6BCF5F70",
x"6D496018",
x"6FBC6135",
x"72FF62B7",
x"76DF6489",
x"7B2B6699",
x"7FB768D6",
x"845A6B30",
x"88FE6D9D",
x"8D907013",
x"9205728C",
x"965774FC",
x"9A857760",
x"9E8779A8",
x"A2577BC9",
x"A5E97DBC",
x"A9327F75",
x"AC2580F1",
x"AEB38232",
x"B0D68338",
x"B285840E",
x"B3C084BC",
x"B485854D",
x"B4DA85C9",
x"B4C68631",
x"B44D8684",
x"B37E86BB",
x"B26186CC",
x"B10A86AC",
x"AF878654",
x"ADF085BF",
x"AC5D84EE",
x"AAE183EC",
x"A99282C3",
x"A8818187",
x"A7B3804C",
x"A7267F20",
x"A6D27E14",
x"A6A27D2C",
x"A6847C6D",
x"A65E7BD3",
x"A61F7B5B",
x"A5BD7B01",
x"A5367ABD",
x"A4917A8F",
x"A3E17A78",
x"A33F7A79",
x"A2C27A95",
x"A27E7ACB",
x"A2817B19",
x"A2CD7B78",
x"A3557BD9",
x"A4047C28",
x"A4B97C53",
x"A5547C47",
x"A5B37BF4",
x"A5BB7B54",
x"A55D7A6A",
x"A49B7943",
x"A38477F7",
x"A23276A5",
x"A0CF7571",
x"9F81747E",
x"9E7473E8",
x"9DC673C3",
x"9D8D7416",
x"9DCC74DB",
x"9E7A75FE",
x"9F837760",
x"A0C278DE",
x"A2177A51",
x"A35A7B9B",
x"A4737C9F",
x"A54A7D4E",
x"A5D97DA8",
x"A6227DB3",
x"A6337D85",
x"A61F7D33",
x"A5FB7CDB",
x"A5DD7C94",
x"A5D47C6D",
x"A5EE7C71",
x"A62E7CA2",
x"A6957CF5",
x"A71E7D60",
x"A7C27DD1",
x"A8777E37",
x"A9387E8A",
x"A9F77EBD",
x"AAAC7ED1",
x"AB4D7ECA",
x"ABD07EAC",
x"AC287E7F",
x"AC4C7E4C",
x"AC337E14",
x"ABDA7DD7",
x"AB437D95",
x"AA767D46",
x"A9807CE8",
x"A8717C75",
x"A7607BEE",
x"A6597B56",
x"A56A7AB3",
x"A4987A0F",
x"A3DD7975",
x"A32C78EB",
x"A2767875",
x"A1A57815",
x"A0A877C1",
x"9F6E7771",
x"9DF37715",
x"9C32769D",
x"9A3275F8",
x"97FA7517",
x"959073F1",
x"92F6727B",
x"902970B4",
x"8D216E9E",
x"89CC6C3F",
x"862169A1",
x"821566D5",
x"7DAD63EF",
x"78FA6107",
x"74215E3D",
x"6F545BAF",
x"6ACF597B",
x"66DB57BD",
x"63B4568F",
x"619055FE",
x"608F560B",
x"60B756B0",
x"61F957DA",
x"642A596D",
x"67115B43",
x"6A685D3B",
x"6DE95F2F",
x"71566101",
x"7480629B",
x"774663F0",
x"799B64FA",
x"7B8165BB",
x"7D09663A",
x"7E456680",
x"7F4C669A",
x"80326690",
x"8101666C",
x"81BF6635",
x"826C65F5",
x"830365B4",
x"837F657A",
x"83DC6553",
x"841B654B",
x"843F656A",
x"845265BA",
x"845D663C",
x"846F66EF",
x"848E67CB",
x"84C468C4",
x"851069C8",
x"85736AC5",
x"85E56BA8",
x"865C6C61",
x"86D26CE5",
x"873B6D2D",
x"87916D3A",
x"87D06D14",
x"87F66CC7",
x"88036C5E",
x"87F96BEB",
x"87DD6B79",
x"87B26B14",
x"877D6AC7",
x"87416A94",
x"86FE6A7F",
x"86BB6A83",
x"86796AA0",
x"86396ACF",
x"86006B0D",
x"85CC6B55",
x"85A06BA1",
x"85796BED",
x"85586C35",
x"853B6C75",
x"851E6CA6",
x"85016CC7",
x"84E36CD5",
x"84C26CCE",
x"84A26CB5",
x"84846C8D",
x"846F6C59",
x"84656C23",
x"846D6BF0",
x"848B6BCB",
x"84C56BB7",
x"851B6BBA",
x"85916BD8",
x"86256C10",
x"86DB6C62",
x"87AE6CCA",
x"88A16D47",
x"89B16DD7",
x"8ADD6E78",
x"8C216F2B",
x"8D746FF0",
x"8ECD70C7",
x"901E71AB",
x"91557297",
x"925D7383",
x"9327745E",
x"939F751A",
x"93BB75A7",
x"937675F5",
x"92D575F6",
x"91E475A9",
x"90BB750C",
x"8F70742A",
x"8E217316",
x"8CE971E5",
x"8BDD70B1",
x"8B0B6F94",
x"8A796EA3",
x"8A1E6DEC",
x"89EF6D76",
x"89DA6D44",
x"89CC6D4A",
x"89B26D7A",
x"89846DC7",
x"893C6E1C",
x"88DD6E68",
x"88726E9E",
x"88036EB8",
x"87A06EB0",
x"87516E85",
x"87186E3B",
x"86F66DDB",
x"86E06D69",
x"86C96CF2",
x"86A76C79",
x"866C6C09",
x"86146BA7",
x"85A16B58",
x"851B6B20",
x"848D6AFF",
x"84046AF5",
x"83876AF9",
x"83176B00",
x"82AA6AFD",
x"822A6ADE",
x"817D6A8F",
x"808169FD",
x"7F1B691D",
x"7D3567E6",
x"7ACB665C",
x"77EB6489",
x"74B56284",
x"715E606A",
x"6E235E5F",
x"6B455C87",
x"69025B04",
x"678759F1",
x"66F05961",
x"6745595D",
x"687659DF",
x"6A625AD7",
x"6CDB5C32",
x"6FAD5DD3",
x"72AA5F9D",
x"75A56173",
x"7883633E",
x"7B2F64EC",
x"7DA46672",
x"7FDF67CC",
x"81E968FA",
x"83C66A02",
x"85816AEB",
x"871A6BBE",
x"88936C83",
x"89EC6D41",
x"8B256DFC",
x"8C3E6EB5",
x"8D3B6F6E",
x"8E1E7021",
x"8EF070CD",
x"8FB77169",
x"907671F0",
x"9131725E",
x"91E272A7",
x"928472CA",
x"930D72BE",
x"93707286",
x"93A47220",
x"939F7192",
x"936270E4",
x"92F07024",
x"92556F65",
x"91A26EB7",
x"90F06E31",
x"90536DE5",
x"8FE66DE2",
x"8FBC6E33",
x"8FE36EDB",
x"90646FD7",
x"9143711A",
x"927B7293",
x"9407742F",
x"95D675D2",
x"97DD776B",
x"9A0B78E5",
x"9C4D7A37",
x"9E927B58",
x"A0C87C49",
x"A2DD7D0C",
x"A4C27DAD",
x"A66A7E36",
x"A7CD7EB0",
x"A8E77F23",
x"A9BC7F99",
x"AA518011",
x"AAB5808B",
x"AAF88108",
x"AB2F8185",
x"AB6D8200",
x"ABC58278",
x"AC4782F1",
x"AD048370",
x"AE0783FA",
x"AF5B8498",
x"B1088550",
x"B3148627",
x"B57E871F",
x"B8458833",
x"BB60895F",
x"BEBF8A93",
x"C2448BC2",
x"C5CE8CD9",
x"C9328DC8",
x"CC408E83",
x"CECB8EFE",
x"D0AD8F3C",
x"D1CA8F3E",
x"D2158F0E",
x"D1928EBC",
x"D05A8E59",
x"CE8F8DF4",
x"CC628D9A",
x"CA058D4E",
x"C7A68D14",
x"C56F8CE6",
x"C3818CBB",
x"C1EA8C88",
x"C0B08C45",
x"BFD08BEA",
x"BF418B79",
x"BEF58AF3",
x"BEDE8A66",
x"BEED89DA",
x"BF16895D",
x"BF4B88FA",
x"BF7E88B4",
x"BF9C8887",
x"BF92886C",
x"BF4B8850",
x"BEAF8824",
x"BDAC87D4",
x"BC368750",
x"BA4C868F",
x"B7F5858F",
x"B54A8457",
x"B26A82F7",
x"AF7D8180",
x"ACAD8008",
x"AA1B7EA3",
x"A7E17D5B",
x"A6087C36",
x"A4817B26",
x"A32E7A1D",
x"A1D978FB",
x"A045779F",
x"9E2C75E8",
x"9B5673BA",
x"97927105",
x"92CF6DCA",
x"8D146A19",
x"868B6617",
x"7F8061F6",
x"784F5DF4",
x"71665A53",
x"6B345750",
x"661C551E",
x"626853DE",
x"604853A1",
x"5FC5545D",
x"60C855F4",
x"631E583C",
x"667D5AF7",
x"6A915DEA",
x"6F0460D5",
x"73876384",
x"77DD65CF",
x"7BD9679E",
x"7F5F68E6",
x"826669B4",
x"84F36A1D",
x"87146A41",
x"88DC6A47",
x"8A646A54",
x"8BC26A8C",
x"8D0A6B04",
x"8E536BCF",
x"8FAB6CEE",
x"91216E55",
x"92B96FF2",
x"947971AB",
x"96567362",
x"984674FE",
x"9A347664",
x"9C077786",
x"9DA5785E",
x"9EFA78EA",
x"9FF17934",
x"A0847947",
x"A0B57936",
x"A091790B",
x"A02978D6",
x"9F9B78A0",
x"9EFE786F",
x"9E6A7846",
x"9DF07826",
x"9D97780F",
x"9D5F7801",
x"9D4277F9",
x"9D3177FC",
x"9D217805",
x"9D077813",
x"9CDA7825",
x"9C9B7833",
x"9C497839",
x"9BED782F",
x"9B8E780D",
x"9B3477D4",
x"9AE07782",
x"9A95771B",
x"9A5576A9",
x"9A177637",
x"99D975D1",
x"99947583",
x"99487555",
x"98F3754A",
x"98957560",
x"9832758D",
x"97CD75C6",
x"976975FC",
x"97017620",
x"96947626",
x"961C7606",
x"959575BD",
x"94F7754D",
x"944074BB",
x"93767412",
x"929D735E",
x"91C672A9",
x"910471FE",
x"906D7166",
x"901770E9",
x"9015708C",
x"90797054",
x"91437043",
x"9274705E",
x"93FD70A7",
x"95C3711F",
x"97AB71C4",
x"99917290",
x"9B50737E",
x"9CC7747B",
x"9DDD7579",
x"9E807667",
x"9EA97730",
x"9E6077CA",
x"9DB6782A",
x"9CC77851",
x"9BB97844",
x"9AB17815",
x"99D577D5",
x"9949779D",
x"99287783",
x"9983779B",
x"9A5A77EB",
x"9BA67878",
x"9D56793D",
x"9F497A2C",
x"A15F7B30",
x"A3737C39",
x"A5647D33",
x"A7177E11",
x"A8777ECA",
x"A97B7F5D",
x"AA257FCF",
x"AA7B8026",
x"AA91806D",
x"AA7480A8",
x"AA3680DA",
x"A9E48101",
x"A9808114",
x"A9058107",
x"A86380C9",
x"A77F8049",
x"A6407F78",
x"A4817E49",
x"A2297CB4",
x"9F227AB9",
x"9B667861",
x"96FB75BA",
x"920172DA",
x"8CA06FDB",
x"870E6CDE",
x"81936A02",
x"7C6D6768",
x"77E0652A",
x"7420635F",
x"71536215",
x"6F8D6155",
x"6ECE6117",
x"6F066155",
x"701661F9",
x"71D262ED",
x"74106418",
x"76A36563",
x"796066B8",
x"7C2A6804",
x"7EE9693E",
x"818E6A5F",
x"84146B69",
x"86796C62",
x"88C16D54",
x"8AEF6E47",
x"8D076F47",
x"8F0A7057",
x"90F47179",
x"92C072AA",
x"946573DF",
x"95D37508",
x"96FE7612",
x"97D976EA",
x"9859777E",
x"987A77C0",
x"983C77AD",
x"97A9774A",
x"96D776A2",
x"95E275CE",
x"94E774EB",
x"940D7419",
x"93767378",
x"933E7321",
x"93767326",
x"94227389",
x"95397444",
x"96A57540",
x"98467664",
x"99FA778F",
x"9BA278A5",
x"9D27798E",
x"9E7E7A3C",
x"9FAF7AB2",
x"A0CA7AF9",
x"A1ED7B2C",
x"A3367B64",
x"A4C57BBF",
x"A6A87C54",
x"A8E37D35",
x"AB667E61",
x"AE0D7FD0",
x"B0AE816D",
x"B3118318",
x"B50784B1",
x"B6648615",
x"B716872C",
x"B71887E4",
x"B67F8839",
x"B5748835",
x"B42987E7",
x"B2D9876E",
x"B1BC86E7",
x"B101866E",
x"B0C98621",
x"B1238614",
x"B20E8652",
x"B37A86DE",
x"B54A87B9",
x"B75D88D4",
x"B98E8A24",
x"BBB98B94",
x"BDC28D10",
x"BF8E8E83",
x"C10B8FDB",
x"C22C9106",
x"C2ED91F4",
x"C34A929D",
x"C34792F9",
x"C2EE9309",
x"C24792CE",
x"C1619253",
x"C04991A5",
x"BF0B90CF",
x"BDB38FDF",
x"BC448EDC",
x"BAC38DCF",
x"B92B8CB6",
x"B7728B90",
x"B5988A58",
x"B3948905",
x"B16B8799",
x"AF2C8615",
x"ACED8484",
x"AACD82F8",
x"A8F48188",
x"A78F8051",
x"A6C37F6D",
x"A6AE7EF1",
x"A7597EEA",
x"A8BF7F54",
x"AAC28025",
x"AD2E8140",
x"AFC68280",
x"B23F83BC",
x"B45484CA",
x"B5C48588",
x"B66785E0",
x"B62585C8",
x"B5048543",
x"B3218468",
x"B0A98353",
x"ADD98221",
x"AAEA80F0",
x"A80D7FD3",
x"A5607ED3",
x"A2ED7DEA",
x"A0A17D02",
x"9E547C01",
x"9BCC7AC1",
x"98CA7922",
x"95127708",
x"907D7467",
x"8AFA7144",
x"849E6DB7",
x"7D9D69E8",
x"764B6607",
x"6F106252",
x"68625F03",
x"62AE5C48",
x"5E525A46",
x"5B8F5911",
x"5A8258A6",
x"5B1F58F5",
x"5D3859DD",
x"60875B35",
x"64AE5CD0",
x"69515E8A",
x"6E10603E",
x"72A361D9",
x"76CF634E",
x"7A76649B",
x"7D8665C6",
x"800466D8",
x"81FE67D3",
x"838468BF",
x"84AB6999",
x"85846A58",
x"861B6AF5",
x"867E6B62",
x"86B76B99",
x"86D16B97",
x"86DC6B63",
x"86EA6B09",
x"870B6A9C",
x"87536A35",
x"87CB69ED",
x"887969D9",
x"89566A03",
x"8A536A6D",
x"8B596B10",
x"8C496BD8",
x"8D016CAD",
x"8D666D72",
x"8D636E0C",
x"8CEF6E69",
x"8C106E7F",
x"8AD66E51",
x"89626DE9",
x"87D96D5F",
x"86666CCD",
x"852F6C4B",
x"84536BEF",
x"83E96BC7",
x"83F36BD7",
x"846C6C14",
x"853E6C72",
x"86486CD7",
x"87666D2D",
x"88736D5B",
x"894F6D52",
x"89E06D0D",
x"8A1B6C8D",
x"89FE6BE1",
x"89956B1C",
x"88F26A58",
x"882E69AE",
x"87666937",
x"86AF6901",
x"861E6916",
x"85BB696F",
x"85846A00",
x"85736AB8",
x"85776B79",
x"85836C28",
x"85806CAD",
x"85636CEF",
x"85246CE3",
x"84BE6C86",
x"84386BDE",
x"839A6AF9",
x"82F469F2",
x"825368E1",
x"81C567E3",
x"81566713",
x"810A6683",
x"80E5663F",
x"80E36649",
x"80FD669A",
x"812A6720",
x"815D67C9",
x"818D687D",
x"81AF6927",
x"81BC69B5",
x"81AD6A1A",
x"817D6A4F",
x"812B6A56",
x"80B96A31",
x"802B69EB",
x"7F89698A",
x"7EDB691D",
x"7E2D68AA",
x"7D8E6838",
x"7D0B67CE",
x"7CB26770",
x"7C906724",
x"7CAD66EC",
x"7D0E66CB",
x"7DB766C5",
x"7EA166DE",
x"7FC56716",
x"8117676C",
x"828667DF",
x"84006868",
x"857368FD",
x"86CC6994",
x"87FC6A20",
x"88F46A97",
x"89AD6AEF",
x"8A1F6B21",
x"8A4B6B2A",
x"8A2F6B09",
x"89D26AC4",
x"89376A5F",
x"886069E1",
x"87516952",
x"860468B8",
x"84776814",
x"82A46766",
x"808166AD",
x"7E0B65E0",
x"7B4164FA",
x"782763F4",
x"74D162CC",
x"7156617E",
x"6DDF6015",
x"6A935E9A",
x"67A45D21",
x"65415BBF",
x"638D5A8D",
x"62A859A2",
x"629D5915",
x"636958F0",
x"64F65939",
x"672359ED",
x"69C05AFB",
x"6C9B5C4F",
x"6F835DCF",
x"724B5F5D",
x"74D160E2",
x"76FF6248",
x"78CC6383",
x"7A3D648B",
x"7B5C6568",
x"7C416621",
x"7CFF66C2",
x"7DAB675B",
x"7E5867F6",
x"7F0E689D",
x"7FD56952",
x"80A86A10",
x"81836AD1",
x"825C6B89",
x"832B6C2D",
x"83E76CB4",
x"848B6D19",
x"85186D59",
x"85906D7A",
x"85FD6D83",
x"866C6D80",
x"86EA6D7C",
x"87866D86",
x"884C6DA4",
x"89456DE1",
x"8A736E3B",
x"8BCF6EB4",
x"8D506F44",
x"8EE46FE2",
x"90767086",
x"91F17126",
x"933F71B4",
x"944F722B",
x"95127288",
x"958372C4",
x"95A272E2",
x"957972E4",
x"951172CD",
x"947E72A4",
x"93D37270",
x"9322723A",
x"927B7206",
x"91F071DA",
x"918871BD",
x"914971B0",
x"913471B7",
x"914371CF",
x"916F71F5",
x"91AB7223",
x"91E97250",
x"921B726E",
x"92327274",
x"92277257",
x"91F1720F",
x"9195719A",
x"911A70FE",
x"908A7044",
x"8FFA6F7F",
x"8F7C6EC7",
x"8F226E35",
x"8F006DE3",
x"8F1B6DE5",
x"8F7A6E47",
x"90176F0D",
x"90E4702A",
x"91D3718D",
x"92CF7316",
x"93C274A5",
x"949E7616",
x"9557774B",
x"95E77832",
x"964F78BC",
x"969478EE",
x"96C178D1",
x"96DC787C",
x"96F47809",
x"970D778F",
x"972C7726",
x"975376DE",
x"978076BE",
x"97AC76C4",
x"97D676E8",
x"97F7771D",
x"980B7751",
x"98117777",
x"9804777F",
x"97E67762",
x"97B3771F",
x"976D76B4",
x"970E762A",
x"9697758C",
x"960774E5",
x"955D7440",
x"949C73AA",
x"93CC732D",
x"92EF72CE",
x"92117290",
x"91387276",
x"9070727E",
x"8FBF729F",
x"8F2972D2",
x"8EAE7310",
x"8E4B734B",
x"8DF4737B",
x"8DA07390",
x"8D3C7382",
x"8CB87345",
x"8BFD72D0",
x"8AFA7217",
x"899B7116",
x"87D56FC7",
x"859E6E27",
x"82F66C38",
x"7FE76A03",
x"7C846797",
x"78EB650A",
x"75426277",
x"71BB6003",
x"6E875DD3",
x"6BDB5C0D",
x"69E35AD3",
x"68C45A3D",
x"68935A59",
x"69545B25",
x"6AF65C8E",
x"6D5C5E76",
x"705560B1",
x"73AB630E",
x"7721655E",
x"7A806772",
x"7D9A6927",
x"80496A6D",
x"82816B3E",
x"843F6BA7",
x"85936BBF",
x"86986BAA",
x"87726B89",
x"88426B7F",
x"892D6BAA",
x"8A486C1A",
x"8BA26CD8",
x"8D3F6DDE",
x"8F116F1E",
x"91047086",
x"92FB71FB",
x"94D77365",
x"967874AD",
x"97C675C6",
x"98AE769F",
x"99277736",
x"99357789",
x"98E677A0",
x"98537782",
x"979A773A",
x"96DA76D5",
x"96357660",
x"95C875E5",
x"95A7756F",
x"95DF7506",
x"967374B3",
x"97587476",
x"987B7457",
x"99C37451",
x"9B147464",
x"9C4C748B",
x"9D5274C1",
x"9E0D74FF",
x"9E71753D",
x"9E7A7572",
x"9E317599",
x"9DA475AA",
x"9CEA75A5",
x"9C1F7588",
x"9B607555",
x"9AC37516",
x"9A5F74D0",
x"9A397490",
x"9A567462",
x"9AAE744E",
x"9B2F745B",
x"9BC6748C",
x"9C5A74DE",
x"9CD67548",
x"9D2475C0",
x"9D3B7633",
x"9D177693",
x"9CBC76D4",
x"9C3676E8",
x"9B9A76D0",
x"9AFD768C",
x"9A747625",
x"9A1275A7",
x"99E47525",
x"99ED74A9",
x"9A287440",
x"9A8773F1",
x"9AF473BE",
x"9B5973A3",
x"9B987396",
x"9B9E7390",
x"9B597389",
x"9AC27376",
x"99DD7358",
x"98B9732D",
x"976A72F8",
x"960B72BE",
x"94B87285",
x"938B7250",
x"9297721C",
x"91E771E8",
x"917E71B1",
x"91557170",
x"91637123",
x"919870C8",
x"91EC7069",
x"9252700D",
x"92C96FC5",
x"93526FA4",
x"93F16FB9",
x"94AF7012",
x"959470B7",
x"96A271A9",
x"97D672DB",
x"9924743B",
x"9A7A75B0",
x"9BC2771B",
x"9CE0785B",
x"9DB97957",
x"9E3B79F8",
x"9E577A32",
x"9E0B7A02",
x"9D5D7971",
x"9C5F788D",
x"9B21776F",
x"99BE7630",
x"984974E8",
x"96CD73AF",
x"95537290",
x"93D07196",
x"923670BB",
x"906E6FF5",
x"8E626F33",
x"8BFD6E62",
x"89346D6F",
x"86096C4A",
x"828D6AEC",
x"7EE06959",
x"7B2F679B",
x"77B165C8",
x"749A63FD",
x"721A6258",
x"705660F7",
x"6F635FF4",
x"6F455F64",
x"6FEC5F4C",
x"713C5FAC",
x"73106079",
x"753E61A2",
x"779E6310",
x"7A1064AE",
x"7C7D6665",
x"7EDD6824",
x"812E69DF",
x"83796B8F",
x"85CC6D31",
x"88356EC5",
x"8AC47051",
x"8D8071D5",
x"906A7358",
x"938074DA",
x"96B67658",
x"99FA77D4",
x"9D367946",
x"A0547AA6",
x"A33F7BEF",
x"A5E07D18",
x"A82B7E19",
x"AA157EF0",
x"ABA17F94",
x"ACD2800C",
x"ADB6805B",
x"AE66808C",
x"AEF480AC",
x"AF7B80C9",
x"B00E80F4",
x"B0BF813D",
x"B19481B2",
x"B28C8256",
x"B3A2832B",
x"B4C48429",
x"B5E18542",
x"B6E18660",
x"B7B7876E",
x"B8568856",
x"B8BD8904",
x"B8F2896A",
x"B9058987",
x"B908895C",
x"B91588FA",
x"B93F8876",
x"B99987E9",
x"BA29876C",
x"BAF08718",
x"BBE186FD",
x"BCE58721",
x"BDE3877E",
x"BEB68808",
x"BF3D88A5",
x"BF5B8938",
x"BEFA89A4",
x"BE0B89CA",
x"BC8F899D",
x"BA93890E",
x"B8328824",
x"B58E86F1",
x"B2D68592",
x"B03D842B",
x"ADF782E7",
x"AC3381EA",
x"AB198154",
x"AAC3813C",
x"AB3B81A6",
x"AC78828A",
x"AE6083CF",
x"B0CC8550",
x"B37F86E4",
x"B63F885C",
x"B8C6898E",
x"BADD8A5A",
x"BC548AA8",
x"BD0C8A71",
x"BCFB89BE",
x"BC2688A2",
x"BAAB873F",
x"B8AF85B9",
x"B6608438",
x"B3EE82DD",
x"B18481C2",
x"AF4280F4",
x"AD3F8075",
x"AB81803D",
x"AA028033",
x"A8B9803F",
x"A7948040",
x"A681801E",
x"A5747FC0",
x"A4647F1C",
x"A3507E32",
x"A23C7D06",
x"A12F7BB0",
x"A0337A46",
x"9F5278E4",
x"9E8A77A2",
x"9DDC7696",
x"9D3F75CB",
x"9CA77546",
x"9C0474FF",
x"9B4974EB",
x"9A6D74F8",
x"996F750F",
x"98527520",
x"9722751A",
x"95F474F5",
x"94DC74AD",
x"93ED7446",
x"933473C3",
x"92B47330",
x"92637292",
x"922971EE",
x"91E77140",
x"916F7082",
x"90956FA7",
x"8F316EA0",
x"8D246D5F",
x"8A606BD8",
x"86EA6A04",
x"82DE67E9",
x"7E666593",
x"79BF6318",
x"752E609D",
x"70F75E43",
x"6D585C32",
x"6A825A8B",
x"6893596A",
x"679658E0",
x"678258F0",
x"683E5992",
x"69A35AB2",
x"6B865C31",
x"6DB85DEC",
x"70105FC1",
x"726D6190",
x"74B7633E",
x"76DC64BA",
x"78D965FC",
x"7AAB6706",
x"7C5967E0",
x"7DE66899",
x"7F58693F",
x"80B169E1",
x"81F46A8C",
x"83246B44",
x"843C6C0C",
x"85416CDE",
x"86326DB3",
x"87116E7C",
x"87E56F2E",
x"88AE6FBB",
x"8973701D",
x"8A35704B",
x"8AF67048",
x"8BB47019",
x"8C6C6FC5",
x"8D156F5C",
x"8DAE6EEE",
x"8E2A6E88",
x"8E876E38",
x"8EC16E0A",
x"8ED76E05",
x"8ECC6E26",
x"8EA56E6B",
x"8E696ECB",
x"8E226F3A",
x"8DDB6FAD",
x"8D9A7014",
x"8D637065",
x"8D3E7099",
x"8D2770AA",
x"8D1D7099",
x"8D1A7069",
x"8D187024",
x"8D126FD1",
x"8D046F7E",
x"8CED6F31",
x"8CCC6EF6",
x"8CA26ED2",
x"8C796EC8",
x"8C506ED5",
x"8C2E6EF9",
x"8C146F2A",
x"8C036F64",
x"8BF76F9A",
x"8BEC6FC8",
x"8BDC6FE6",
x"8BC06FF0",
x"8B9A6FE8",
x"8B696FCB",
x"8B316FA3",
x"8AF96F73",
x"8ACB6F43",
x"8AB16F1A",
x"8AB16EFF",
x"8AD06EF3",
x"8B0D6EF6",
x"8B5F6F06",
x"8BBC6F1C",
x"8C146F30",
x"8C586F3A",
x"8C746F31",
x"8C606F13",
x"8C116EDB",
x"8B876E8A",
x"8AC66E26",
x"89D66DB5",
x"88C86D44",
x"87A86CD9",
x"868A6C82",
x"85806C42",
x"84956C21",
x"83D66C20",
x"83496C38",
x"82F36C65",
x"82CE6C9C",
x"82D56CD4",
x"82FA6CFF",
x"83316D13",
x"83696D08",
x"83916CD7",
x"83976C7C",
x"83726BF6",
x"83176B49",
x"82846A7A",
x"81B96991",
x"80C16897",
x"7FA26796",
x"7E6F669B",
x"7D3165B1",
x"7BF764E0",
x"7ACF6434",
x"79BE63AB",
x"78CB634B",
x"77F6630D",
x"773F62ED",
x"76A462E2",
x"761E62E0",
x"75AA62DD",
x"753B62CC",
x"74C962A4",
x"74486259",
x"73A761E9",
x"72D96149",
x"71CB607C",
x"70705F7C",
x"6EBF5E4B",
x"6CB45CED",
x"6A585B67",
x"67BD59C7",
x"64FA5819",
x"62375670",
x"5F9C54E3",
x"5D525387",
x"5B805275",
x"5A4451BF",
x"59B15172",
x"59CA5195",
x"5A855222",
x"5BCB5309",
x"5D7D5439",
x"5F785591",
x"619456F7",
x"63B2584F",
x"65BA5982",
x"67975A87",
x"69425B59",
x"6ABA5BFD",
x"6C005C7E",
x"6D1D5CF1",
x"6E165D62",
x"6EEC5DDD",
x"6FA45E69",
x"703B5F03",
x"70AD5F9F",
x"70F76031",
x"711960A4",
x"711060EA",
x"70E260F7",
x"709660C6",
x"7035605C",
x"6FCC5FC6",
x"6F685F1A",
x"6F135E6C",
x"6ED55DD6",
x"6EB45D6E",
x"6EB15D41",
x"6ECC5D56",
x"6F025DAB",
x"6F4B5E35",
x"6FA15EE7",
x"6FFF5FAB",
x"705C606E",
x"70B5611F",
x"710761B1",
x"7151621A",
x"71906259",
x"71C86272",
x"71FA626A",
x"7228624F",
x"7253622B",
x"72806207",
x"72B061EC",
x"72E261DF",
x"731861E2",
x"735261F3",
x"7390620E",
x"73D2622D",
x"741A6248",
x"7466625C",
x"74BA6266",
x"75146262",
x"75776250",
x"75DF6234",
x"764A620D",
x"76B061DF",
x"770B61AD",
x"77556179",
x"77846143",
x"77946110",
x"777F60DF",
x"774560B5",
x"76ED6097",
x"7681608B",
x"760F609D",
x"75A460D2",
x"75546134",
x"752B61C5",
x"75376289",
x"757D6376",
x"76006483",
x"76BB659E",
x"77A166B5",
x"78A867B4",
x"79C16886",
x"7ADC691E",
x"7BEF6977",
x"7CED6994",
x"7DD3697D",
x"7E9E6947",
x"7F4E6904",
x"7FE068CC",
x"805868B2",
x"80B568C4",
x"80F76904",
x"811B696F",
x"812169F7",
x"810A6A89",
x"80D96B10",
x"80966B78",
x"804C6BB1",
x"800C6BB7",
x"7FE36B8D",
x"7FE36B3E",
x"801A6AE1",
x"80906A8C",
x"81456A56",
x"82346A51",
x"834E6A89",
x"847C6AFA",
x"85A86B9C",
x"86B56C57",
x"878E6D12",
x"88206DB4",
x"88636E24",
x"88596E55",
x"880D6E3F",
x"87916DE9",
x"86FD6D62",
x"86666CBE",
x"85DD6C13",
x"856C6B72",
x"850B6AE5",
x"84AC6A6C",
x"843269F9",
x"8376697A",
x"825368D6",
x"80A867F5",
x"7E5F66BF",
x"7B73652E",
x"77F66345",
x"740D6115",
x"6FED5EBD",
x"6BDE5C61",
x"68235A2C",
x"65025846",
x"62AD56CD",
x"614555DA",
x"60D25574",
x"61415599",
x"626C563A",
x"64195740",
x"660A588F",
x"68055A0A",
x"69D45B94",
x"6B535D14",
x"6C765E7A",
x"6D3D5FB7",
x"6DBB60BF",
x"6E106191",
x"6E5C6229",
x"6EBE628D",
x"6F4F62BF",
x"701B62C8",
x"712162B1",
x"72586286",
x"73AB6253",
x"75036227",
x"764A620D",
x"77696213",
x"7855623C",
x"79096291",
x"7983630D",
x"79CB63AB",
x"79E96462",
x"79EA6523",
x"79D965E0",
x"79BA668D",
x"7996671A",
x"796D6780",
x"794567B8",
x"792167C5",
x"790367AB",
x"78F06775",
x"78F0672B",
x"790C66DF",
x"7947669B",
x"79A7666A",
x"7A2F6656",
x"7AE06660",
x"7BB7668A",
x"7CAB66D2",
x"7DB56731",
x"7ECC67A3",
x"7FE36823",
x"80F268A8",
x"81ED6932",
x"82CE69BA",
x"83906A3E",
x"842E6AB8",
x"84AA6B26",
x"85036B82",
x"85416BCA",
x"856A6BF9",
x"85896C10",
x"85A76C0F",
x"85CF6BFD",
x"860B6BE3",
x"865F6BCF",
x"86CF6BCB",
x"87586BE3",
x"87F46C23",
x"889D6C8C",
x"89486D1C",
x"89EA6DCA",
x"8A7E6E88",
x"8B016F45",
x"8B736FF2",
x"8BD8707F",
x"8C3970E5",
x"8C9E7120",
x"8D0E7134",
x"8D90712E",
x"8E22711A",
x"8EC17108",
x"8F637102",
x"8FFD7110",
x"90807137",
x"90DF716F",
x"911171AF",
x"911071E9",
x"90DA7210",
x"90797219",
x"8FF071FB",
x"8F4C71B5",
x"8E9B714B",
x"8DE670C5",
x"8D387030",
x"8C956F97",
x"8C076F09",
x"8B8D6E90",
x"8B2B6E31",
x"8AE76DF3",
x"8AC56DD7",
x"8ACB6DD8",
x"8AFD6DF6",
x"8B636E2D",
x"8BFA6E75",
x"8CBC6EC8",
x"8D9E6F1E",
x"8E8A6F6E",
x"8F676FAE",
x"901A6FD5",
x"90866FD9",
x"90936FB7",
x"90376F6E",
x"8F6D6F02",
x"8E456E80",
x"8CD36DF8",
x"8B386D7C",
x"89976D1A",
x"880E6CE2",
x"86B46CD4",
x"858E6CE9",
x"84976D12",
x"83B26D31",
x"82B86D27",
x"817C6CD2",
x"7FCE6C16",
x"7D896ADF",
x"7A966928",
x"76F366FC",
x"72BB6474",
x"6E1761B7",
x"69485EEE",
x"64975C4D",
x"604E59FE",
x"5CB35824",
x"59F656D7",
x"583D5622",
x"578A55FE",
x"57D25660",
x"58F2572C",
x"5AB85849",
x"5CEF5995",
x"5F5F5AF6",
x"61D45C50",
x"64265D90",
x"663A5EA7",
x"68025F8B",
x"69776039",
x"6AA360B2",
x"6B8E60FD",
x"6C4C611F",
x"6CE96127",
x"6D75611D",
x"6DFC610E",
x"6E866101",
x"6F1760FC",
x"6FB260FE",
x"70556108",
x"70FC6114",
x"71A16117",
x"723D610A",
x"72C760E7",
x"733860AE",
x"738D6060",
x"73C16004",
x"73D85FA9",
x"73D65F5C",
x"73C85F2E",
x"73BB5F2C",
x"73BF5F63",
x"73E55FD5",
x"7437607D",
x"74BB6153",
x"75756248",
x"765B6345",
x"77606437",
x"78726507",
x"797965A5",
x"7A606607",
x"7B166628",
x"7B8D660A",
x"7BC265BB",
x"7BB56548",
x"7B7264C6",
x"7B096449",
x"7A8C63E5",
x"7A0E63A5",
x"79A26395",
x"795663B4",
x"793163FD",
x"79356463",
x"795F64D9",
x"79A8654E",
x"7A0365AF",
x"7A6665F3",
x"7AC46611",
x"7B146609",
x"7B4E65DE",
x"7B70659D",
x"7B7A6550",
x"7B736509",
x"7B6064D3",
x"7B4F64BB",
x"7B4B64C8",
x"7B5E64FD",
x"7B946558",
x"7BF365D3",
x"7C7F6669",
x"7D31670E",
x"7E0467BA",
x"7EEB6860",
x"7FD268FA",
x"80AB6980",
x"816669EB",
x"81F76A3A",
x"825A6A6B",
x"82916A80",
x"82A16A7C",
x"82986A62",
x"82846A38",
x"82746A03",
x"827469C8",
x"82876989",
x"82AB6948",
x"82D96907",
x"830368C4",
x"8318687D",
x"830B6832",
x"82D367E3",
x"826C6791",
x"81DC673E",
x"813266EF",
x"808066AA",
x"7FDD6675",
x"7F5D6655",
x"7F0E6650",
x"7EF56668",
x"7F0D6699",
x"7F4966DF",
x"7F946732",
x"7FD6678D",
x"7FF767E0",
x"7FE96828",
x"7FA4685C",
x"7F2A6876",
x"7E8A6876",
x"7DD8685B",
x"7D2B6826",
x"7C9567D6",
x"7C24676C",
x"7BD866E5",
x"7BA5663F",
x"7B746579",
x"7B28648D",
x"7AA36380",
x"79C56256",
x"7883611D",
x"76DC5FE3",
x"74E65EC3",
x"72C45DD3",
x"70A85D2C",
x"6ECF5CE4",
x"6D705D06",
x"6CBA5D95",
x"6CCF5E8B",
x"6DB85FD9",
x"6F706164",
x"71D86314",
x"74C564CC",
x"78076679",
x"7B6F680C",
x"7ED2697F",
x"82176ADB",
x"85346C2A",
x"882A6D7D",
x"8B0D6EE6",
x"8DF17073",
x"90F4722A",
x"942B740C",
x"979F7615",
x"9B567834",
x"9F427A60",
x"A34F7C85",
x"A7607E9B",
x"AB568095",
x"AF0E8276",
x"B26E843B",
x"B56185E6",
x"B7DB877A",
x"B9D688F6",
x"BB578A55",
x"BC6D8B8E",
x"BD2A8C9B",
x"BDAA8D6F",
x"BE0C8E03",
x"BE6E8E58",
x"BEF58E73",
x"BFC08E63",
x"C0E78E41",
x"C27E8E24",
x"C4898E2A",
x"C7018E6A",
x"C9D38EF6",
x"CCDB8FD3",
x"CFEF90FE",
x"D2E29266",
x"D58893F3",
x"D7BA958A",
x"D964970C",
x"DA829864",
x"DB209982",
x"DB629A5E",
x"DB749AFF",
x"DB859B6E",
x"DBC79BBA",
x"DC629BF6",
x"DD6B9C2D",
x"DEE19C68",
x"E0B09CA4",
x"E2B19CDB",
x"E4AC9CFF",
x"E6659CFD",
x"E79F9CC7",
x"E8279C4B",
x"E7DE9B85",
x"E6B89A75",
x"E4C19926",
x"E21D97AA",
x"DF01961D",
x"DBB0949A",
x"D8759342",
x"D592922E",
x"D3479176",
x"D1BA9125",
x"D1039142",
x"D12091C4",
x"D1F7929A",
x"D35893AB",
x"D50B94D9",
x"D6C89602",
x"D8509700",
x"D96297B8",
x"D9D39811",
x"D98697FC",
x"D8729772",
x"D6A29676",
x"D4309514",
x"D143935E",
x"CE069168",
x"CAA38F4B",
x"C73F8D1B",
x"C3F48AEC",
x"C0D388CC",
x"BDE486C5",
x"BB2284DC",
x"B8858315",
x"B6078171",
x"B39E7FF2",
x"B1497E99",
x"AF0C7D68",
x"ACF37C64",
x"AB087B92",
x"A95F7AF7",
x"A8087A96",
x"A7127A74",
x"A6837A8C",
x"A6567ADE",
x"A6817B5D",
x"A6ED7BFB",
x"A77B7CAA",
x"A8087D54",
x"A8707DE4",
x"A88E7E47",
x"A84C7E70",
x"A7997E51",
x"A67A7DEB",
x"A4FA7D44",
x"A3397C67",
x"A1597B67",
x"9F817A5A",
x"9DD27950",
x"9C607857",
x"9B2E7775",
x"9A2B76A3",
x"992F75D1",
x"980774E4",
x"967673BD",
x"943F723D",
x"9135704A",
x"8D3F6DD8",
x"88666AE8",
x"82CE678D",
x"7CBB63F2",
x"768A604B",
x"70A35CD7",
x"6B6F59DA",
x"674B578F",
x"647D5625",
x"632A55B8",
x"6352564C",
x"64D557CF",
x"67755A18",
x"6AE25CEE",
x"6EBE6011",
x"72B1633E",
x"766F6634",
x"79B868C5",
x"7C686ACC",
x"7E6C6C3E",
x"7FCC6D17",
x"80986D6B",
x"80F26D51",
x"80F96CEB",
x"80D16C58",
x"809B6BB7",
x"80726B20",
x"80666AA1",
x"80876A48",
x"80D66A17",
x"81566A0F",
x"82016A2B",
x"82CC6A69",
x"83AE6AC2",
x"849A6B31",
x"85816BAE",
x"86596C30",
x"87176CAD",
x"87B46D19",
x"882A6D66",
x"88796D8A",
x"88A56D7D",
x"88B56D3D",
x"88AF6CCA",
x"889E6C2D",
x"88886B76",
x"88796ABA",
x"88736A10",
x"887E698D",
x"889D6947",
x"88D0694B",
x"891B69A0",
x"897D6A42",
x"89F46B2A",
x"8A806C45",
x"8B1E6D7D",
x"8BCB6EBA",
x"8C816FE4",
x"8D3E70E5",
x"8DF971AF",
x"8EAE7237",
x"8F56727B",
x"8FEE727F",
x"9071724D",
x"90DD71F0",
x"912E7176",
x"916270EF",
x"91797066",
x"91736FE5",
x"91506F72",
x"91136F10",
x"90BC6EBF",
x"90566E7D",
x"8FE66E48",
x"8F776E1D",
x"8F126DFA",
x"8EC26DE1",
x"8E906DCF",
x"8E816DCB",
x"8E956DD2",
x"8EC86DE9",
x"8F106E0C",
x"8F606E3A",
x"8FAB6E6C",
x"8FE26E9E",
x"8FFA6ECD",
x"8FEE6EF0",
x"8FBE6F0A",
x"8F726F19",
x"8F146F23",
x"8EB56F2D",
x"8E666F43",
x"8E316F69",
x"8E1E6FAD",
x"8E31700F",
x"8E627092",
x"8EA77131",
x"8EF471E6",
x"8F3B72A4",
x"8F727361",
x"8F92740D",
x"8F9F74A0",
x"8FA17510",
x"8FA7755B",
x"8FBF7582",
x"8FFC7586",
x"90637571",
x"90FB7548",
x"91BB7516",
x"929474DC",
x"937074A0",
x"94367461",
x"94D0741A",
x"952973CB",
x"9538736F",
x"94FD7302",
x"947E7282",
x"93CD71F4",
x"92FA715A",
x"921870BA",
x"912F701A",
x"90456F7E",
x"8F506EE8",
x"8E436E54",
x"8D086DBA",
x"8B8A6D12",
x"89B96C51",
x"87916B6B",
x"85186A5E",
x"82656928",
x"7F9A67D5",
x"7CE56675",
x"7A74651D",
x"787363E8",
x"770662ED",
x"76416246",
x"762561FC",
x"76AB6214",
x"77B86289",
x"792A6349",
x"7AE06444",
x"7CBB6563",
x"7EA56696",
x"809467CC",
x"82866904",
x"84876A3F",
x"86A56B86",
x"88F46CE6",
x"8B806E68",
x"8E557013",
x"917171E8",
x"94CF73DF",
x"985D75EA",
x"9C0777F2",
x"9FB579E5",
x"A34F7BAF",
x"A6C07D40",
x"A9F67E91",
x"ACE47FA3",
x"AF848080",
x"B1D68132",
x"B3DD81C9",
x"B5A08256",
x"B72982E3",
x"B882837A",
x"B9BA841F",
x"BADA84D4",
x"BBF18598",
x"BD078669",
x"BE228745",
x"BF49882C",
x"C07B891D",
x"C1B28A14",
x"C2E48B0D",
x"C4048C01",
x"C5018CE5",
x"C5C68DA8",
x"C6468E3C",
x"C6708E93",
x"C6408EA1",
x"C5B68E63",
x"C4DE8DDB",
x"C3D08D14",
x"C2A88C24",
x"C18F8B25",
x"C0AB8A35",
x"C025896D",
x"C01988E7",
x"C09D88B2",
x"C1B588D4",
x"C34C894C",
x"C5468A0A",
x"C7718AFA",
x"C9968C06",
x"CB788D10",
x"CCE48E03",
x"CDAF8EC8",
x"CDC38F53",
x"CD228F9E",
x"CBE48FAB",
x"CA368F84",
x"C8568F35",
x"C6848ED2",
x"C5028E6D",
x"C4058E17",
x"C3B28DDC",
x"C4128DC3",
x"C5198DD2",
x"C6A58E00",
x"C8848E49",
x"CA788EA1",
x"CC498EFE",
x"CDC18F59",
x"CEC18FAA",
x"CF368FF0",
x"CF22902D",
x"CE959065",
x"CDAF909D",
x"CC9090D5",
x"CB5B910D",
x"CA26913F",
x"C8FE9163",
x"C7E5916A",
x"C6D19148",
x"C5B390F2",
x"C478905D",
x"C3128F8E",
x"C17B8E8A",
x"BFB78D5D",
x"BDD38C1D",
x"BBE58ADA",
x"BA0F89AC",
x"B86A889F",
x"B70F87BF",
x"B6148708",
x"B57E8678",
x"B5498603",
x"B5688597",
x"B5C68525",
x"B64684A5",
x"B6CA840E",
x"B73A8361",
x"B77F82A3",
x"B78881E0",
x"B74C8123",
x"B6CA8078",
x"B6087FEA",
x"B50C7F7B",
x"B3E67F2B",
x"B29E7EF1",
x"B13B7EBD",
x"AFBD7E7E",
x"AE1F7E1E",
x"AC507D87",
x"AA337CA5",
x"A7A67B64",
x"A48779B9",
x"A0B2779F",
x"9C117515",
x"969B7226",
x"905D6EE6",
x"897C6B72",
x"823167E9",
x"7ACF6474",
x"73B4613B",
x"6D3D5E62",
x"67C45C08",
x"63925A45",
x"60D45922",
x"5F96589C",
x"5FC858A8",
x"613A592C",
x"63A75A0B",
x"66BB5B24",
x"6A215C57",
x"6D8A5D8B",
x"70B55EAE",
x"73795FB5",
x"75BC609F",
x"777D6177",
x"78C76243",
x"79AF6313",
x"7A5363EF",
x"7ACC64E0",
x"7B3165E6",
x"7B9166FA",
x"7BF96814",
x"7C6A6923",
x"7CEC6A14",
x"7D7C6ADB",
x"7E1B6B6C",
x"7ECB6BBE",
x"7F8C6BD4",
x"805C6BB1",
x"813B6B63",
x"82206AF9",
x"83046A86",
x"83DC6A19",
x"849869C1",
x"852C698A",
x"858D6977",
x"85B56989",
x"85A469BA",
x"855D6A02",
x"84F06A54",
x"846D6AA7",
x"83E76AF0",
x"83746B2A",
x"83276B4F",
x"830B6B62",
x"832A6B63",
x"83846B5E",
x"84136B57",
x"84C96B58",
x"85986B69",
x"86706B90",
x"87416BD1",
x"87FD6C2A",
x"889E6C99",
x"89216D19",
x"89886DA0",
x"89D86E26",
x"8A156E9E",
x"8A486F00",
x"8A706F43",
x"8A916F5F",
x"8AA56F55",
x"8AA76F24",
x"8A936ED4",
x"8A666E6C",
x"8A246DF9",
x"89D56D8C",
x"89886D31",
x"89556CF6",
x"89526CE6",
x"89986D08",
x"8A376D59",
x"8B366DDB",
x"8C946E85",
x"8E3E6F4A",
x"9018701F",
x"91FD70F6",
x"93C271C3",
x"953F7279",
x"96557312",
x"96EA7385",
x"96F873CD",
x"968773E8",
x"95A573D7",
x"94737399",
x"930D7334",
x"919572AA",
x"90257203",
x"8ECF7144",
x"8D9C7075",
x"8C8A6FA0",
x"8B8E6ECA",
x"8A9D6DFD",
x"89A56D3E",
x"889E6C92",
x"87816BFC",
x"86506B7D",
x"85156B16",
x"83E36AC8",
x"82CE6A94",
x"81EF6A7A",
x"81596A7C",
x"811D6A9C",
x"81426ADB",
x"81C66B38",
x"829B6BB2",
x"83AB6C44",
x"84D66CDF",
x"85FC6D7C",
x"86F96E08",
x"87B46E75",
x"88156EB4",
x"88176EBD",
x"87B76E89",
x"87046E17",
x"86106D70",
x"84F36CA0",
x"83C26BB2",
x"828B6AB8",
x"815869BA",
x"801D68BF",
x"7ECB67C5",
x"7D4566C6",
x"7B6C65B5",
x"79246481",
x"76586321",
x"73066188",
x"6F3B5FB8",
x"6B1E5DBC",
x"66E65BA8",
x"62DB599C",
x"5F4A57BD",
x"5C7F5633",
x"5ABA5521",
x"5A2754A3",
x"5AD854CD",
x"5CC255A1",
x"5FC25712",
x"639C590C",
x"68055B6D",
x"6CAE5E0D",
x"714F60C1",
x"75A86363",
x"798D65D2",
x"7CE667F5",
x"7FAF69BC",
x"81F76B24",
x"83D66C2E",
x"856A6CE3",
x"86CD6D55",
x"88186D93",
x"89566DB0",
x"8A8B6DBD",
x"8BAE6DC7",
x"8CB16DD7",
x"8D846DF0",
x"8E1A6E16",
x"8E696E41",
x"8E6D6E69",
x"8E2C6E86",
x"8DB66E92",
x"8D1E6E83",
x"8C796E59",
x"8BDC6E17",
x"8B596DC1",
x"8AFB6D61",
x"8AC56D00",
x"8AB16CA8",
x"8AB16C62",
x"8AAF6C2D",
x"8A936C09",
x"8A456BF0",
x"89AE6BDB",
x"88BE6BBF",
x"87706B97",
x"85C86B5B",
x"83D66B0D",
x"81B46AB2",
x"7F816A52",
x"7D6569F9",
x"7B8069B2",
x"79F66987",
x"78DD697F",
x"7845699C",
x"783069DC",
x"78906A38",
x"79526AA7",
x"7A586B1D",
x"7B7C6B8D",
x"7C9D6BED",
x"7D9B6C35",
x"7E5F6C61",
x"7ED96C6D",
x"7F076C5B",
x"7EF36C30",
x"7EAC6BF2",
x"7E4C6BA8",
x"7DE86B5C",
x"7D956B14",
x"7D626AD4",
x"7D526A9E",
x"7D606A73",
x"7D7D6A4E",
x"7D946A28",
x"7D9469FF",
x"7D6C69CC",
x"7D176991",
x"7C9E6954",
x"7C1B691E",
x"7BB46901",
x"7B966910",
x"7BF06961",
x"7CED6A04",
x"7EAC6B04",
x"81356C62",
x"847C6E13",
x"885A7005",
x"8C9E7219",
x"9108742F",
x"95577623",
x"995077DA",
x"9CC7793E",
x"9FA27A4A",
x"A1DA7AFE",
x"A37A7B64",
x"A4977B93",
x"A54C7B9C",
x"A5B17B92",
x"A5D67B81",
x"A5C67B6B",
x"A57E7B50",
x"A4F77B25",
x"A4267ADE",
x"A30B7A75",
x"A1A879E4",
x"A00A792D",
x"9E4D785E",
x"9C947785",
x"9B0376B9",
x"99BE760C",
x"98E07592",
x"987A7554",
x"988D7552",
x"99057588",
x"99CA75E4",
x"9AB57652",
x"9B9A76BD",
x"9C507710",
x"9CB3773A",
x"9CA2772C",
x"9C0876DE",
x"9AD3764B",
x"98FE7572",
x"96887451",
x"937972EA",
x"8FDD713E",
x"8BCE6F55",
x"87696D34",
x"82D66AEB",
x"7E446886",
x"79E86620",
x"75F363D0",
x"729A61B5",
x"70035FE6",
x"6E4A5E7C",
x"6D785D83",
x"6D865D02",
x"6E595CF8",
x"6FCC5D57",
x"71AE5E0D",
x"73CC5F00",
x"75F9601A",
x"780D6143",
x"79EF6268",
x"7B91637C",
x"7CF66477",
x"7E28655B",
x"7F386625",
x"803966E0",
x"813C6791",
x"824C683C",
x"836C68EB",
x"849A699C",
x"85CE6A52",
x"86FA6B0F",
x"88136BCC",
x"89086C8A",
x"89D66D42",
x"8A766DF0",
x"8AE66E8F",
x"8B2C6F14",
x"8B506F7C",
x"8B5C6FC0",
x"8B596FD9",
x"8B556FC7",
x"8B536F89",
x"8B5D6F24",
x"8B746E9E",
x"8B986E05",
x"8BC46D62",
x"8BF16CC7",
x"8C186C41",
x"8C316BDE",
x"8C346BA7",
x"8C1D6B9E",
x"8BE76BC4",
x"8B986C10",
x"8B346C76",
x"8AC46CE3",
x"8A526D48",
x"89EA6D90",
x"899A6DAD",
x"89696D97",
x"895F6D4D",
x"897D6CD2",
x"89C36C3A",
x"8A2F6B96",
x"8AB86AFF",
x"8B586A8F",
x"8C066A59",
x"8CBE6A6F",
x"8D7A6AD9",
x"8E366B97",
x"8EF06C9D",
x"8FA76DD9",
x"90596F37",
x"9107709D",
x"91B171F6",
x"92567330",
x"92FA743D",
x"939B7519",
x"943C75C3",
x"94DF763E",
x"95817693",
x"962576C7",
x"96C876E1",
x"976276E4",
x"97ED76D0",
x"986276A3",
x"98B4765D",
x"98D975F8",
x"98CA7579",
x"988574E1",
x"98077434",
x"9753737F",
x"967472C8",
x"9576721D",
x"94637186",
x"934C710A",
x"923C70AE",
x"91397070",
x"904C704E",
x"8F737041",
x"8EAF7041",
x"8DFE7045",
x"8D5C7043",
x"8CC97034",
x"8C457014",
x"8BD36FDE",
x"8B796F92",
x"8B386F33",
x"8B146EC5",
x"8B0B6E4F",
x"8B186DD9",
x"8B346D6C",
x"8B4C6D0F",
x"8B536CC5",
x"8B356C94",
x"8AE36C7C",
x"8A556C75",
x"89866C7A",
x"887A6C82",
x"87426C7F",
x"85F16C68",
x"84A16C37",
x"836A6BE5",
x"82606B72",
x"81916ADE",
x"80FC6A30",
x"8097696B",
x"80466897",
x"7FEC67B7",
x"7F5C66CB",
x"7E7265D2",
x"7D0B64CB",
x"7B1463B1",
x"788A6280",
x"757C613C",
x"72105FEA",
x"6E795E95",
x"6AF75D4C",
x"67CF5C21",
x"653F5B26",
x"637C5A73",
x"62A65A11",
x"62CA5A0D",
x"63DB5A66",
x"65B85B17",
x"68335C12",
x"6B105D48",
x"6E145EA1",
x"710A6008",
x"73C96169",
x"763862B1",
x"784E63D5",
x"7A1164D0",
x"7B9665A0",
x"7CF46649",
x"7E4B66D8",
x"7FAC6756",
x"812A67D3",
x"82C4685C",
x"847768FC",
x"863269BA",
x"87E56A9A",
x"89796B9A",
x"8ADC6CB1",
x"8C066DD4",
x"8CEF6EF3",
x"8D9C6FFC",
x"8E1870DF",
x"8E6F718D",
x"8EAC7200",
x"8EE07230",
x"8F117220",
x"8F4571D8",
x"8F7C7161",
x"8FB570CE",
x"8FED702D",
x"901F6F92",
x"904B6F0C",
x"906E6EA9",
x"908E6E72",
x"90AE6E6F",
x"90D06E9E",
x"90FA6EFE",
x"912E6F80",
x"916A701C",
x"91AF70BE",
x"91F47158",
x"923571D7",
x"92697230",
x"928B7258",
x"9294724B",
x"9281720D",
x"924F71A6",
x"92007123",
x"91947092",
x"910E7005",
x"90766F86",
x"8FCF6F21",
x"8F226ED8",
x"8E776EAA",
x"8DD76E90",
x"8D496E82",
x"8CD96E73",
x"8C8B6E5F",
x"8C666E3E",
x"8C6A6E0F",
x"8C986DD7",
x"8CEA6D9C",
x"8D5B6D69",
x"8DE06D47",
x"8E716D3E",
x"8F076D54",
x"8F9B6D88",
x"90276DD7",
x"90A86E38",
x"911E6EA1",
x"91856F03",
x"91DF6F52",
x"92276F83",
x"92596F90",
x"92716F75",
x"926A6F35",
x"92426ED8",
x"91F46E68",
x"91856DF8",
x"90FD6D94",
x"90666D51",
x"8FCD6D3A",
x"8F466D58",
x"8EDC6DAD",
x"8E9D6E37",
x"8E8D6EEB",
x"8EAC6FB7",
x"8EF1708A",
x"8F4F714E",
x"8FB271F0",
x"900D7262",
x"904D729A",
x"9069729A",
x"905F7268",
x"902F720F",
x"8FE771A3",
x"8F927133",
x"8F3F70D1",
x"8EFC7088",
x"8ED2705C",
x"8EC6704F",
x"8ED9705C",
x"8F077076",
x"8F4B7094",
x"8F9D70AB",
x"8FF470B5",
x"904C70AD",
x"909D7094",
x"90DF706C",
x"9104703A",
x"90FE6FFC",
x"90B86FB4",
x"90146F59",
x"8EF76EE2",
x"8D466E3B",
x"8AE76D54",
x"87D26C1E",
x"84096A8F",
x"7F9E68A4",
x"7AB86666",
x"758D63EC",
x"705C6152",
x"6B6F5EBF",
x"67075C5C",
x"63635A4D",
x"60AE58B5",
x"5F0357A8",
x"5E69572E",
x"5ED45740",
x"602657D1",
x"623458C6",
x"64CF5A00",
x"67C55B61",
x"6AE65CCF",
x"6E065E32",
x"71045F7E",
x"73C760AB",
x"763B61BB",
x"785C62AE",
x"7A25638A",
x"7B9B6455",
x"7CC86513",
x"7DB865C6",
x"7E7D6670",
x"7F2B6710",
x"7FDB67AA",
x"809E683F",
x"818E68D6",
x"82B86975",
x"84276A20",
x"85DB6ADE",
x"87CB6BB0",
x"89E36C92",
x"8C076D7F",
x"8E146E69",
x"8FE96F43",
x"915F6FFE",
x"925D708C",
x"92D070E2",
x"92B470FC",
x"920E70DA",
x"90F67082",
x"8F877000",
x"8DE76F62",
x"8C3E6EB7",
x"8AAC6E0A",
x"894F6D69",
x"88396CD8",
x"87706C5B",
x"86EF6BF2",
x"86AA6B9A",
x"868A6B52",
x"867C6B17",
x"86696AE9",
x"86416AC8",
x"85F76AB5",
x"858A6AB5",
x"84FF6AC7",
x"84626AEC",
x"83C16B26",
x"832E6B6D",
x"82BC6BC1",
x"82796C19",
x"826D6C6F",
x"829E6CBB",
x"830A6CF9",
x"83AB6D27",
x"84766D41",
x"855D6D4D",
x"86536D4D",
x"874B6D47",
x"883B6D45",
x"891A6D51",
x"89E96D70",
x"8AA76DAA",
x"8B596E02",
x"8C096E7A",
x"8CBC6F12",
x"8D7E6FC1",
x"8E567085",
x"8F467152",
x"90527220",
x"917372E8",
x"92A273A1",
x"93D37447",
x"94FA74D4",
x"96047548",
x"96E375A3",
x"978875E2",
x"97EC7606",
x"9804760F",
x"97D075F8",
x"975375BE",
x"96917561",
x"959474DE",
x"94697437",
x"931D7372",
x"91BC7297",
x"905971B7",
x"8F0170E2",
x"8DC2702B",
x"8CAB6FA7",
x"8BC56F64",
x"8B1D6F6C",
x"8AB56FC4",
x"8A907065",
x"8AAB713E",
x"8AFD723D",
x"8B797344",
x"8C0D7436",
x"8CA574F6",
x"8D2F756F",
x"8D98758F",
x"8DD0754D",
x"8DD274AD",
x"8D9573B9",
x"8D217285",
x"8C797126",
x"8BA76FB5",
x"8AB46E4D",
x"89A76CF9",
x"887E6BC8",
x"873B6ABE",
x"85D269D6",
x"84376903",
x"825C6838",
x"80376762",
x"7DC26670",
x"7B006555",
x"77FD640A",
x"74CE628D",
x"719160E6",
x"6E695F24",
x"6B7C5D59",
x"68EC5B9E",
x"66D55A08",
x"654958AF",
x"645157A4",
x"63E656F1",
x"63F9569C",
x"647056A5",
x"653156FF",
x"661D57A1",
x"671A5878",
x"68135973",
x"68FC5A81",
x"69CF5B92",
x"6A8F5C9C",
x"6B445D95",
x"6BF85E7A",
x"6CB35F46",
x"6D7C5FFC",
x"6E586098",
x"6F41611F",
x"70316191",
x"711A61EF",
x"71F06235",
x"72A76268",
x"73356286",
x"73946291",
x"73C76290",
x"73D26287",
x"73C56280",
x"73AF6281",
x"73A36295",
x"73B162C1",
x"73E6630A",
x"744F636D",
x"74EC63E9",
x"75B86473",
x"76A864FD",
x"77AA6577",
x"78A765D2",
x"798965FF",
x"7A3865F2",
x"7AA365A7",
x"7AC16521",
x"7A8C646C",
x"7A0C6397",
x"794E62B7",
x"786B61E3",
x"7779612F",
x"769360AE",
x"75D16066",
x"7544605C",
x"74F46086",
x"74E260D6",
x"75026138",
x"75456198",
x"759661E0",
x"75DE6203",
x"760A61F9",
x"761061C3",
x"75E6616C",
x"75916101",
x"751A609B",
x"7490604D",
x"7404602B",
x"738A6041",
x"732E6091",
x"72F7611B",
x"72EC61D0",
x"7304629F",
x"733A6372",
x"73826431",
x"73CF64CB",
x"741B6532",
x"745F6560",
x"7499655B",
x"74CB652A",
x"74FF64DE",
x"75386489",
x"7581643B",
x"75DE6404",
x"764F63EC",
x"76CF63F4",
x"7756641D",
x"77D66458",
x"783F649E",
x"788164DF",
x"7891650E",
x"78666525",
x"77FC651E",
x"775964F9",
x"768A64B7",
x"759D6460",
x"74AA63FA",
x"73C4638D",
x"72FF631E",
x"726B62B2",
x"720E6248",
x"71ED61E2",
x"7200617E",
x"723E611F",
x"729460C3",
x"72F5606E",
x"734C6024",
x"73915FE6",
x"73BA5FB9",
x"73BF5F9F",
x"73A55F97",
x"736F5F9A",
x"73215F9F",
x"72C25F9F",
x"72595F8E",
x"71EB5F64",
x"71755F18",
x"70F95EAB",
x"70755E1E",
x"6FE35D7B",
x"6F415CCC",
x"6E865C1E",
x"6DAD5B7A",
x"6CB05AE9",
x"6B895A6E",
x"6A315A05",
x"68A459A8",
x"66E05949",
x"64E958DD",
x"62C75857",
x"608757B3",
x"5E4456F0",
x"5C175614",
x"5A21552C",
x"5886544A",
x"57645382",
x"56D152E8",
x"56DF528C",
x"57905278",
x"58DB52B3",
x"5AA95336",
x"5CDC53FB",
x"5F5254F1",
x"61E35608",
x"646D572C",
x"66D4584C",
x"68FC5957",
x"6ADB5A43",
x"6C665B07",
x"6DA05B9E",
x"6E8C5C08",
x"6F315C4C",
x"6F9A5C6E",
x"6FD45C7B",
x"6FE65C7E",
x"6FE05C87",
x"6FCF5C9F",
x"6FBE5CD5",
x"6FB85D2C",
x"6FC65DA9",
x"6FF25E4C",
x"703C5F08",
x"70A65FD8",
x"712A60A8",
x"71BF616D",
x"725F6218",
x"72FF629F",
x"739362FC",
x"7416632E",
x"74846338",
x"74DF6321",
x"752A62F6",
x"756862BE",
x"759B6284",
x"75CB6253",
x"75F56232",
x"76166222",
x"762A6227",
x"762D6241",
x"7619626D",
x"75EC62AB",
x"75A862F4",
x"75556348",
x"74FD639D",
x"74B263F2",
x"7486643E",
x"7489647F",
x"74C964AE",
x"755264CB",
x"762164D2",
x"772E64C5",
x"786664A5",
x"79AF6474",
x"7AED6437",
x"7BFF63ED",
x"7CC6639A",
x"7D316341",
x"7D3162E2",
x"7CC56280",
x"7BFA621E",
x"7AE861BF",
x"79AB6168",
x"7869611D",
x"774660E6",
x"766560C9",
x"75D860C9",
x"75B160E7",
x"75EC6127",
x"76806180",
x"775861F2",
x"78536272",
x"795362F9",
x"7A39637D",
x"7AEC63FA",
x"7B586469",
x"7B7664C6",
x"7B486511",
x"7ADC6548",
x"7A44656C",
x"7996657D",
x"78E7657C",
x"784C6569",
x"77D56541",
x"77836504",
x"775864B1",
x"774B6449",
x"774E63CC",
x"77526341",
x"774B62AD",
x"772B6218",
x"76EF6193",
x"76996124",
x"762E60D9",
x"75BF60BB",
x"755E60CE",
x"75196115",
x"7502618E",
x"75236232",
x"758162F4",
x"761A63C8",
x"76DF649B",
x"77C16562",
x"78A86609",
x"797C6687",
x"7A2366D3",
x"7A8966E9",
x"7AA166C6",
x"7A65666F",
x"79D565E9",
x"78F9653E",
x"77DF6477",
x"7699639E",
x"753462BE",
x"73C161DD",
x"72496106",
x"70D5603B",
x"6F635F80",
x"6DF55ED6",
x"6C895E3F",
x"6B205DB9",
x"69C15D45",
x"68785CE1",
x"67565C92",
x"66725C59",
x"65E35C39",
x"65BF5C38",
x"66145C5C",
x"66E95CA7",
x"68375D1B",
x"69EF5DBB",
x"6BF85E81",
x"6E315F69",
x"707C606C",
x"72BB617E",
x"74DE6298",
x"76DE63B2",
x"78C264C6",
x"7AA065D8",
x"7C9366E6",
x"7EBE67FD",
x"813C6926",
x"84256A6B",
x"87806BD4",
x"8B466D69",
x"8F5D6F2A",
x"93A1710F",
x"97E0730B",
x"9BE9750B",
x"9F8B76FC",
x"A29F78C8",
x"A50E7A5E",
x"A6D07BAF",
x"A7EE7CB4",
x"A8807D74",
x"A8A47DF2",
x"A87E7E43",
x"A8337E74",
x"A7E17E9B",
x"A79E7EC6",
x"A7717EFC",
x"A75D7F45",
x"A75A7F9E",
x"A75D7FFC",
x"A757805A",
x"A74280A8",
x"A71580DD",
x"A6D680F2",
x"A68A80E7",
x"A63F80BD",
x"A605807E",
x"A5EB8032",
x"A5FB7FE7",
x"A63D7FA8",
x"A6B07F7E",
x"A74F7F6E",
x"A80B7F78",
x"A8D77F9B",
x"A99F7FCD",
x"AA518002",
x"AADD802D",
x"AB368042",
x"AB4F802D",
x"AB227FE8",
x"AAAC7F6A",
x"A9ED7EB0",
x"A8EA7DBC",
x"A7A87C98",
x"A6307B51",
x"A48F79FF",
x"A2D578B4",
x"A10E7786",
x"9F497689",
x"9D9775C8",
x"9C01754B",
x"9A91750F",
x"99497509",
x"982B7527",
x"97337557",
x"965D7585",
x"95A4759D",
x"95017596",
x"9473756A",
x"93F9751D",
x"939574BB",
x"934C7452",
x"932273F5",
x"931B73B3",
x"9338739A",
x"937773B1",
x"93D373F9",
x"9443746C",
x"94BB74FF",
x"953175A2",
x"95987648",
x"95EA76E4",
x"9622776C",
x"964377DA",
x"9650782D",
x"96527868",
x"9652788D",
x"965C78A3",
x"967A78AC",
x"96B378AA",
x"970B789C",
x"9783787F",
x"98157851",
x"98BC780F",
x"996977B4",
x"9A107746",
x"9A9B76C6",
x"9AFB763C",
x"9B1F75B1",
x"9AF7752F",
x"9A7974BD",
x"999F745F",
x"986E741A",
x"96F373EA",
x"953C73C6",
x"936573A3",
x"91837379",
x"8FAE7337",
x"8DF672D2",
x"8C607240",
x"8AE37176",
x"896C706F",
x"87D96F24",
x"86036D93",
x"83C26BBB",
x"80F2699D",
x"7D7D673C",
x"796064A3",
x"74AF61DA",
x"6F945EF7",
x"6A4E5C11",
x"65275946",
x"607356B8",
x"5C835485",
x"599752D0",
x"57DF51AF",
x"57715133",
x"58415160",
x"5A31522D",
x"5D095388",
x"60825550",
x"64515761",
x"682A5992",
x"6BCC5BBD",
x"6F075DBF",
x"71BB5F7E",
x"73DC60EC",
x"75706201",
x"768B62C4",
x"774C633F",
x"77D26386",
x"784163AB",
x"78B263C1",
x"793F63D6",
x"79EF63F7",
x"7AC7642A",
x"7BBC646C",
x"7CC564BC",
x"7DCE6513",
x"7EC16566",
x"7F9165B1",
x"802F65ED",
x"8097661A",
x"80CB663B",
x"80D26658",
x"80BB6679",
x"809A66AA",
x"807E66F5",
x"8076675C",
x"808C67E5",
x"80BE6889",
x"8107693F",
x"815969F9",
x"81A16AA4",
x"81CE6B2D",
x"81CF6B84",
x"819A6B9E",
x"812E6B76",
x"80936B0F",
x"7FD66A73",
x"7F1169B4",
x"7E5C68E9",
x"7DCF682B",
x"7D83678E",
x"7D816728",
x"7DD26703",
x"7E706720",
x"7F4E677D",
x"8058680D",
x"817768BF",
x"82976982",
x"839F6A41",
x"84816AF0",
x"85316B84",
x"85AB6BFA",
x"85EF6C54",
x"86006C97",
x"85E66CCA",
x"85AE6CF3",
x"855D6D19",
x"85016D3B",
x"84A26D58",
x"84466D6B",
x"83F46D6E",
x"83B26D59",
x"83816D2B",
x"83656CE3",
x"83586C84",
x"83596C17",
x"83626BA4",
x"836D6B37",
x"83736AD9",
x"836C6A90",
x"83536A5E",
x"83276A42",
x"82E46A37",
x"82906A32",
x"822E6A2D",
x"81C56A1D",
x"815C69FD",
x"80F969C9",
x"809D6983",
x"8049692E",
x"7FFA68CC",
x"7FA86868",
x"7F4C6801",
x"7EDC67A0",
x"7E506742",
x"7DAA66E8",
x"7CE6668E",
x"7C0D6635",
x"7B2765D8",
x"7A426576",
x"79686511",
x"78A664AB",
x"77FF644B",
x"777963F4",
x"770E63AB",
x"76B76376",
x"766A6353",
x"761E6344",
x"75C66342",
x"755F634B",
x"74E66352",
x"745F6355",
x"73CF6349",
x"733F632A",
x"72B562F0",
x"723A629B",
x"71CB6225",
x"7165618E",
x"70FD60D3",
x"70865FF4",
x"6FED5EF1",
x"6F215DC8",
x"6E115C7A",
x"6CB05B0D",
x"6AF65984",
x"68E657EB",
x"6687564F",
x"63EC54BF",
x"612B534A",
x"5E635205",
x"5BBA50FC",
x"59525040",
x"574F4FD7",
x"55D14FC4",
x"54EE5009",
x"54B3509D",
x"55215175",
x"56305282",
x"57C553B5",
x"59C054FA",
x"5BFB5643",
x"5E4A577F",
x"608558A5",
x"628D59AB",
x"644B5A8D",
x"65B35B47",
x"66C75BDF",
x"67935C59",
x"682A5CBD",
x"68A65D15",
x"691E5D6A",
x"69A75DC3",
x"6A4F5E29",
x"6B1D5E9D",
x"6C0A5F1B",
x"6D0E5FA1",
x"6E1A6024",
x"6F1B609B",
x"700360FC",
x"70C5613E",
x"715C615F",
x"71C76160",
x"720D614B",
x"723E6128",
x"72666108",
x"729860FE",
x"72E56117",
x"7355615A",
x"73ED61CE",
x"74AF6269",
x"75936321",
x"768D63E5",
x"778C649E",
x"7881653B",
x"796065AD",
x"7A2065EA",
x"7ABB65F5",
x"7B3865D6",
x"7B9D65A0",
x"7BFA6565",
x"7C5F6538",
x"7CDC652E",
x"7D7C654F",
x"7E45659D",
x"7F356614",
x"803F66A5",
x"81536741",
x"825667D2",
x"832F6848",
x"83C46896",
x"840168B5",
x"83DF68A8",
x"835D6876",
x"828A682B",
x"817E67D5",
x"805B6781",
x"7F46673C",
x"7E66670D",
x"7DDC66F7",
x"7DC166F9",
x"7E1D670E",
x"7EEF6732",
x"8027675F",
x"81AA678E",
x"835267BC",
x"84F967EB",
x"867A6814",
x"87B5683E",
x"88936869",
x"89046894",
x"890D68C2",
x"88B268F2",
x"88086923",
x"87246954",
x"86206983",
x"851469B2",
x"841369DE",
x"832E6A06",
x"826F6A28",
x"81D86A44",
x"81696A55",
x"811E6A5B",
x"80F06A51",
x"80D66A37",
x"80C86A0A",
x"80BE69CC",
x"80B2697D",
x"80A16923",
x"808668BE",
x"80636858",
x"803867F5",
x"80096799",
x"7FD56746",
x"7F9E6703",
x"7F6766CC",
x"7F2E66A0",
x"7EF0667D",
x"7EAB6662",
x"7E586648",
x"7DF56631",
x"7D7D661A",
x"7CEF6600",
x"7C4C65E5",
x"7B9665C5",
x"7ACE659E",
x"79F96570",
x"791A6534",
x"783064E8",
x"77386486",
x"762E640A",
x"75096376",
x"73BF62C6",
x"724B6200",
x"70A86129",
x"6EDB6048",
x"6CEC5F63",
x"6AED5E87",
x"68FB5DB8",
x"67305CFE",
x"65AD5C60",
x"648D5BE0",
x"63E85B81",
x"63CB5B45",
x"64355B2C",
x"651E5B39",
x"66705B6B",
x"68105BC5",
x"69DC5C43",
x"6BB45CE6",
x"6D7D5DA7",
x"6F215E80",
x"70995F69",
x"71DD6056",
x"72FC613E",
x"73FC6215",
x"74EF62D6",
x"75E26379",
x"76E06400",
x"77F2646D",
x"791664C8",
x"7A49651B",
x"7B836572",
x"7CBB65D2",
x"7DE86642",
x"7F0066C5",
x"80006756",
x"80E267F2",
x"81A4688A",
x"82466917",
x"82C96990",
x"832E69EC",
x"83776A2B",
x"83A86A54",
x"83C96A6C",
x"83E56A87",
x"84096AB1",
x"84456AFD",
x"84AB6B75",
x"854B6C1D",
x"862F6CF5",
x"875C6DEE",
x"88CC6EF6",
x"8A706FF9",
x"8C3470DC",
x"8DFA718C",
x"8FA171F6",
x"91107216",
x"922E71EF",
x"92ED718D",
x"934B7106",
x"93507073",
x"930B6FEB",
x"92946F85",
x"92016F4D",
x"91676F48",
x"90D96F75",
x"905D6FC4",
x"8FF77026",
x"8FA47085",
x"8F5970CE",
x"8F1070F4",
x"8EBE70EF",
x"8E5D70C0",
x"8DED706E",
x"8D707008",
x"8CED6F9C",
x"8C6A6F3D",
x"8BF16EF8",
x"8B8B6ED8",
x"8B3C6EE2",
x"8B0A6F13",
x"8AF36F69",
x"8AFB6FD9",
x"8B21705A",
x"8B6570E1",
x"8BC87165",
x"8C4B71E1",
x"8CF07250",
x"8DB672AD",
x"8E9E72F8",
x"8FA17330",
x"90B67354",
x"91D37364",
x"92E6735C",
x"93DF7340",
x"94AA730D",
x"953672C7",
x"9579726C",
x"95697203",
x"9504718D",
x"94507110",
x"93597090",
x"922C700D",
x"90DC6F8A",
x"8F7C6F06",
x"8E1C6E80",
x"8CD36DF9",
x"8BAB6D70",
x"8AB16CE6",
x"89EC6C5F",
x"89606BE1",
x"89136B72",
x"88FE6B19",
x"89246ADC",
x"897A6AC5",
x"89FA6AD2",
x"8A956B04",
x"8B406B59",
x"8BE96BC8",
x"8C816C45",
x"8CFA6CCA",
x"8D4B6D48",
x"8D696DB7",
x"8D556E0D",
x"8D0D6E44",
x"8C916E54",
x"8BE56E3A",
x"8B036DEF",
x"89E46D6F",
x"887C6CB5",
x"86B76BBD",
x"847F6A7F",
x"81BF68F6",
x"7E696723",
x"7A766506",
x"75EC62A4",
x"70DF600B",
x"6B785D4B",
x"65E55A78",
x"606657AF",
x"5B3B550B",
x"56A452A6",
x"52D7509D",
x"50004F04",
x"4E374DEA",
x"4D834D5A",
x"4DDA4D51",
x"4F1F4DCA",
x"51274EB3",
x"53C24FFB",
x"56BB5185",
x"59DB533A",
x"5CF154FD",
x"5FD556B5",
x"6269584F",
x"649C59BB",
x"66655AF0",
x"67CA5BE9",
x"68DB5CA7",
x"69A85D2C",
x"6A4F5D83",
x"6AE35DB2",
x"6B795DC5",
x"6C215DC5",
x"6CDF5DBC",
x"6DB35DB3",
x"6E935DAF",
x"6F755DB8",
x"70465DCF",
x"70FA5DF7",
x"71865E2F",
x"71E25E78",
x"72115ECF",
x"721C5F2E",
x"72105F92",
x"71FD5FF9",
x"71F6605A",
x"720960B5",
x"72446108",
x"72AA6152",
x"733F6195",
x"740061D5",
x"74E36215",
x"75E2625D",
x"76EF62B1",
x"78046315",
x"791A638E",
x"7A2A641B",
x"7B2F64BA",
x"7C286565",
x"7D106614",
x"7DE066C1",
x"7E946760",
x"7F2567EC",
x"7F8D685C",
x"7FC568B1",
x"7FC968E9",
x"7F9A6907",
x"7F3A6910",
x"7EAE690C",
x"7E0068FD",
x"7D3A68E9",
x"7C6868D2",
x"7B9468B5",
x"7AC7688C",
x"7A06684C",
x"795567F2",
x"78B26770",
x"781E66C2",
x"779465E8",
x"770E64E5",
x"768A63C2",
x"7603628B",
x"757A6155",
x"74EF602F",
x"74655F2C",
x"73DF5E5A",
x"73655DC1",
x"72F95D64",
x"72A15D41",
x"72625D4F",
x"723B5D80",
x"722B5DC9",
x"72305E1A",
x"723F5E67",
x"72535EA8",
x"725F5EDA",
x"72585EFD",
x"72375F12",
x"71F25F22",
x"71865F31",
x"70F55F42",
x"70445F5A",
x"6F7D5F77",
x"6EAE5F9A",
x"6DE85FB9",
x"6D3A5FD3",
x"6CB05FE3",
x"6C565FE4",
x"6C335FD9",
x"6C485FC3",
x"6C905FA9",
x"6D065F92",
x"6DA05F86",
x"6E545F8A",
x"6F175FA5",
x"6FE25FD9",
x"70AE6025",
x"71756084",
x"723260ED",
x"72E66159",
x"738C61C1",
x"7423621B",
x"74A56264",
x"7513629B",
x"756862BF",
x"75A062D0",
x"75BA62D5",
x"75AF62CB",
x"758062B2",
x"75256289",
x"74966248",
x"73CB61E4",
x"72B76155",
x"71516090",
x"6F8C5F8E",
x"6D665E4D",
x"6ADF5CD0",
x"68025B21",
x"64E35950",
x"61A65774",
x"5E7255A9",
x"5B795409",
x"58EE52AF",
x"570251B3",
x"55DB5126",
x"55975115",
x"5640517F",
x"57CE5264",
x"5A2B53B9",
x"5D30556B",
x"60A7576A",
x"645C599C",
x"68115BE6",
x"6B935E2C",
x"6EB26055",
x"714E6241",
x"735263DA",
x"74BA650E",
x"758D65CB",
x"75E0660E",
x"75D165D8",
x"75806538",
x"75136442",
x"74AA6313",
x"746061CB",
x"744B608A",
x"746F5F6E",
x"74CE5E91",
x"75595DFD",
x"75FD5DB9",
x"76A35DC1",
x"772E5E08",
x"778C5E7E",
x"77AD5F11",
x"778E5FB3",
x"77326056",
x"76AD60F4",
x"7610618D",
x"757A6222",
x"750262BB",
x"74BF635A",
x"74C16407",
x"750964C2",
x"75946584",
x"76566649",
x"773B6707",
x"783167B0",
x"7925683A",
x"7A0D689B",
x"7AE268CE",
x"7BA868D2",
x"7C6C68AB",
x"7D3A6862",
x"7E246803",
x"7F38679E",
x"807E6746",
x"81F9670E",
x"839E6703",
x"855D6731",
x"872167A0",
x"88CE684C",
x"8A4B6934",
x"8B836A47",
x"8C676B70",
x"8CF66C9E",
x"8D326DB5",
x"8D2B6EA0",
x"8CF46F4D",
x"8CA76FAE",
x"8C566FBE",
x"8C146F80",
x"8BEC6EFA",
x"8BDC6E3E",
x"8BDA6D5C",
x"8BD96C6D",
x"8BC06B84",
x"8B7D6AB5",
x"8AFA6A0D",
x"8A316996",
x"891D6954",
x"87C66944",
x"8643695F",
x"84AA699A",
x"831869E3",
x"81AD6A2D",
x"807E6A69",
x"7FA16A89",
x"7F1A6A86",
x"7EE96A5E",
x"7F036A14",
x"7F5669B2",
x"7FC96945",
x"804568DB",
x"80B26880",
x"80FD6841",
x"8117681E",
x"80F6681A",
x"809A682D",
x"80036849",
x"7F386865",
x"7E486870",
x"7D3E6865",
x"7C27683B",
x"7B1467F3",
x"7A106793",
x"79256723",
x"785C66AD",
x"77B46637",
x"773065C8",
x"76C86560",
x"767564FD",
x"76306498",
x"75EC642E",
x"75A363B5",
x"754E632E",
x"74E66297",
x"746C61F6",
x"73DE6152",
x"733B60AF",
x"72846017",
x"71BB5F88",
x"70D95F04",
x"6FDF5E80",
x"6ECA5DF6",
x"6D965D5C",
x"6C475CAC",
x"6AE25BE6",
x"69705B0B",
x"68025A2B",
x"66A75956",
x"6575589F",
x"6480581E",
x"63DB57E0",
x"639457F1",
x"63B45854",
x"643E5901",
x"652D59E7",
x"66765AF6",
x"680D5C14",
x"69E15D2C",
x"6BDE5E31",
x"6DF55F15",
x"70165FDA",
x"72356086",
x"744C6122",
x"765661BE",
x"78516264",
x"7A3D6325",
x"7C196403",
x"7DE964FF",
x"7FAB660E",
x"815F672A",
x"8301683F",
x"848E693F",
x"86046A1C",
x"87606ACB",
x"88A56B4C",
x"89D86BA3",
x"8B036BDC",
x"8C346C0A",
x"8D7B6C44",
x"8EE96CA0",
x"908D6D35",
x"92716E16",
x"949C6F4A",
x"970B70D2",
x"99B572A7",
x"9C8674BA",
x"9F6A76F2",
x"A2497934",
x"A5087B65",
x"A7957D6E",
x"A9DF7F39",
x"ABDC80B7",
x"AD8B81E3",
x"AEF582BC",
x"B0258345",
x"B12C8385",
x"B219838A",
x"B2FE835C",
x"B3E78307",
x"B4DC8297",
x"B5DE8216",
x"B6ED818F",
x"B7FC810C",
x"B9028098",
x"B9EE803F",
x"BAB28005",
x"BB3F7FF2",
x"BB8C800A",
x"BB998046",
x"BB6A80A3",
x"BB0B8118",
x"BA93819C",
x"BA218225",
x"B9D082B1",
x"B9C3833F",
x"BA1883D4",
x"BAE3847D",
x"BC2D8540",
x"BDF5862B",
x"C02D8740",
x"C2B68884",
x"C56E89E9",
x"C82C8B60",
x"CACA8CD3",
x"CD278E27",
x"CF2F8F45",
x"D0DA901B",
x"D22A90A1",
x"D33090D6",
x"D40290C8",
x"D4B79087",
x"D565902D",
x"D6168FD2",
x"D6CD8F89",
x"D77E8F5D",
x"D8168F58",
x"D8798F6F",
x"D88B8F97",
x"D8308FBF",
x"D75D8FD3",
x"D6098FC6",
x"D4418F8A",
x"D21C8F1B",
x"CFBD8E7D",
x"CD4B8DB9",
x"CAEF8CE0",
x"C8D18C01",
x"C70E8B32",
x"C5B38A83",
x"C4C98A00",
x"C44789B4",
x"C41E89A2",
x"C43389C9",
x"C46D8A22",
x"C4AD8AA1",
x"C4DB8B34",
x"C4DE8BC9",
x"C4A88C4E",
x"C42D8CAE",
x"C36E8CDC",
x"C26A8CCB",
x"C12B8C77",
x"BFB68BDD",
x"BE1B8B05",
x"BC5B89F6",
x"BA7E88B8",
x"B87B8753",
x"B64785D0",
x"B3D0842C",
x"B0F88267",
x"ADA58077",
x"A9BB7E53",
x"A5257BEF",
x"9FDF7948",
x"99F4765E",
x"93877339",
x"8CCD6FEC",
x"860E6C92",
x"7F9B694E",
x"79CC6644",
x"74F2639B",
x"71496174",
x"6F005FEC",
x"6E255F0E",
x"6EAA5EE2",
x"70685F5F",
x"73286074",
x"76A56209",
x"7A9D6400",
x"7ED3663F",
x"831F68AE",
x"87696B38",
x"8BAA6DD2",
x"8FEE7076",
x"944C7326",
x"98DA75E4",
x"9DAB78B3",
x"A2C67B96",
x"A8247E8C",
x"ADAF818B",
x"B34A848A",
x"B8CC8777",
x"BE0C8A43",
x"C2EB8CDD",
x"C7538F38",
x"CB3A914B",
x"CEA59313",
x"D1A29494",
x"D44695D6",
x"D6A796E5",
x"D8D897CC",
x"DAE29896",
x"DCC69948",
x"DE7C99EB",
x"DFFB9A7B",
x"E1339AF8",
x"E2199B5A",
x"E2A79B9D",
x"E2E29BBD",
x"E2D19BB0",
x"E2829B78",
x"E2099B10",
x"E1789A7D",
x"E0DD99C5",
x"E04198EE",
x"DFAE9805",
x"DF269716",
x"DEAD9634",
x"DE46956F",
x"DDF694DB",
x"DDCB9486",
x"DDD0947D",
x"DE0F94C4",
x"DE909559",
x"DF519633",
x"E044973D",
x"E151985C",
x"E2549975",
x"E3259A68",
x"E3999B1A",
x"E38F9B76",
x"E2EC9B72",
x"E1B09B0D",
x"DFE99A52",
x"DDB99958",
x"DB54983A",
x"D8F19719",
x"D6CE9611",
x"D51C9542",
x"D3FC94BD",
x"D37F948A",
x"D39D94AD",
x"D43B9519",
x"D53095B8",
x"D6449678",
x"D7469737",
x"D80597DF",
x"D85D9856",
x"D83C988D",
x"D79D987C",
x"D6939821",
x"D5379787",
x"D3B096C1",
x"D22695E3",
x"D0C3950C",
x"CFA79453",
x"CEEB93D1",
x"CE9B9393",
x"CEB193A3",
x"CF2393F8",
x"CFD79484",
x"D0AD9533",
x"D18695E3",
x"D246967C",
x"D2D496E2",
x"D3239702",
x"D33196D4",
x"D309965F",
x"D2BD95B4",
x"D26894EE",
x"D226942A",
x"D212938A",
x"D23D932A",
x"D2AD931A",
x"D35D9360",
x"D43993F8",
x"D52694C9",
x"D60195BD",
x"D6A696B1",
x"D6FB9785",
x"D6E7981D",
x"D6649869",
x"D575985F",
x"D42397FF",
x"D27F974C",
x"D0989654",
x"CE72951A",
x"CC0C93A4",
x"C95191EF",
x"C6238FED",
x"C25D8D94",
x"BDD48ACD",
x"B86D878F",
x"B21583D2",
x"AAD67F9C",
x"A2D37B05",
x"9A4C7630",
x"9198714F",
x"891F6CA0",
x"8151685E",
x"7A9164C2",
x"753461FC",
x"71706025",
x"6F5E5F49",
x"6EF05F59",
x"6FFC6038",
x"723A61B9",
x"755963A8",
x"78FD65D2",
x"7CD56804",
x"80986A1D",
x"84146BFF",
x"872C6DA1",
x"89D86F03",
x"8C1E702B",
x"8E147127",
x"8FD57203",
x"917672CA",
x"9310737F",
x"94AF7425",
x"965974B9",
x"980A7537",
x"99BC759D",
x"9B6475EC",
x"9CFA762A",
x"9E777661",
x"9FDA769F",
x"A12476F1",
x"A2577765",
x"A37E7803",
x"A49B78CD",
x"A5B179BA",
x"A6BA7AC1",
x"A7B57BCD",
x"A8917CC9",
x"A9427DA0",
x"A9BB7E41",
x"A9F07E9E",
x"A9DA7EB2",
x"A97A7E7B",
x"A8D77E05",
x"A7FE7D5B",
x"A7017C8E",
x"A5F77BAC",
x"A4F47AC9",
x"A40B79EF",
x"A349792F",
x"A2B6788D",
x"A2557812",
x"A21C77BE",
x"A2077793",
x"A207778D",
x"A21177AA",
x"A21A77E4",
x"A218782F",
x"A2077885",
x"A1E378DB",
x"A1AC7929",
x"A1677968",
x"A1187995",
x"A0C679AD",
x"A07B79B4",
x"A03E79B0",
x"A01479A6",
x"A008799F",
x"A01C799F",
x"A05479AA",
x"A0B079C1",
x"A12E79E4",
x"A1C57A0C",
x"A26D7A3C",
x"A3217A6E",
x"A3D67AA9",
x"A48B7AF2",
x"A53D7B58",
x"A5F37BE8",
x"A6B87CB3",
x"A79C7DC6",
x"A8B27F29",
x"AA1180E4",
x"ABCC82F0",
x"ADF08540",
x"B08787C5",
x"B38E8A64",
x"B6F78D08",
x"BAAB8F94",
x"BE8A91F4",
x"C26A9416",
x"C62095E9",
x"C9879769",
x"CC72988C",
x"CEC79951",
x"D06F99B7",
x"D16299BE",
x"D1A3996B",
x"D14098C1",
x"D04E97CB",
x"CEEC9697",
x"CD399535",
x"CB5493BB",
x"C95B923E",
x"C76790D1",
x"C5868F86",
x"C3C08E65",
x"C2158D70",
x"C07C8CA0",
x"BEEE8BE5",
x"BD578B2C",
x"BBAD8A62",
x"B9E68976",
x"B7FC885D",
x"B5F48717",
x"B3D485AB",
x"B1AD842C",
x"AF8C82AF",
x"AD7F8149",
x"AB8E800B",
x"A9B27EFC",
x"A7DD7E16",
x"A5F07D47",
x"A3C37C6D",
x"A12B7B64",
x"9DF77A02",
x"9A047823",
x"953C75AD",
x"8FA2729C",
x"894F6EF8",
x"82796AE2",
x"7B6A668D",
x"74806238",
x"6E195E28",
x"68935A9C",
x"643857CF",
x"613E55E7",
x"5FBB54F7",
x"5FA454F8",
x"60CF55D1",
x"62FF5756",
x"65E2594C",
x"69265B74",
x"6C795D92",
x"6F975F73",
x"725360EE",
x"749061F4",
x"76486280",
x"778962A1",
x"786C6276",
x"79106221",
x"799661CB",
x"7A166195",
x"7AA4619A",
x"7B4561E6",
x"7BF46279",
x"7CA76346",
x"7D486438",
x"7DC66532",
x"7E146617",
x"7E2766CF",
x"7E006749",
x"7DAA6781",
x"7D38677F",
x"7CC46751",
x"7C68670D",
x"7C3F66CF",
x"7C5E66AE",
x"7CCE66BB",
x"7D9066FF",
x"7E986779",
x"7FD36820",
x"812768DE",
x"827669A0",
x"83A46A4F",
x"849D6ADB",
x"85556B34",
x"85CB6B59",
x"86076B4F",
x"861D6B23",
x"861D6AE3",
x"86216AA3",
x"863E6A73",
x"867E6A62",
x"86ED6A79",
x"87886ABE",
x"88486B2E",
x"89216BC4",
x"8A046C78",
x"8AE26D3D",
x"8BB16E08",
x"8C676ECE",
x"8D036F82",
x"8D81701D",
x"8DE57094",
x"8E3270E6",
x"8E6D710C",
x"8E9A7109",
x"8EB970E1",
x"8ED07097",
x"8EDF703A",
x"8EE76FD1",
x"8EEA6F65",
x"8EE96F02",
x"8EE46EAA",
x"8EDD6E61",
x"8ECF6E23",
x"8EB46DEC",
x"8E876DB4",
x"8E3E6D76",
x"8DD06D2E",
x"8D3B6CDC",
x"8C7B6C86",
x"8B976C33",
x"8A9A6BEF",
x"89946BC8",
x"889B6BCB",
x"87C66BFA",
x"872A6C5B",
x"86D26CE3",
x"86C36D88",
x"86FD6E35",
x"876F6ED5",
x"88016F54",
x"889B6F9F",
x"891F6FAB",
x"89776F72",
x"89916EF6",
x"89636E43",
x"88F06D61",
x"88426C65",
x"876A6B61",
x"867D6A63",
x"858E697A",
x"84B168B1",
x"83F0680D",
x"83506791",
x"82D2673B",
x"82706709",
x"822066F5",
x"81D866F9",
x"81916710",
x"81436734",
x"80EF6762",
x"8094679A",
x"803967DC",
x"7FE9682B",
x"7FA5688C",
x"7F796901",
x"7F62698D",
x"7F5F6A2D",
x"7F666AD9",
x"7F696B87",
x"7F516C20",
x"7F076C8D",
x"7E706CB3",
x"7D766C78",
x"7C036BC4",
x"7A0D6A8C",
x"779468CF",
x"74A36699",
x"71526406",
x"6DC5613C",
x"6A285E6D",
x"66AD5BCB",
x"63865985",
x"60DF57C9",
x"5EDF56AF",
x"5DA05644",
x"5D2A5682",
x"5D7C5751",
x"5E885892",
x"60315A18",
x"62585BB9",
x"64D95D4C",
x"678F5EB1",
x"6A565FD5",
x"6D1160B1",
x"6FA36149",
x"71F761AB",
x"73FD61EC",
x"75AA621F",
x"76F3625A",
x"77D962AA",
x"785C6314",
x"7884639B",
x"7862643B",
x"780764E6",
x"778A6594",
x"77076637",
x"769A66C5",
x"76586738",
x"7655678D",
x"769D67C4",
x"773167E0",
x"780A67E5",
x"791A67D6",
x"7A4967BB",
x"7B7F6796",
x"7CA06768",
x"7D946732",
x"7E4C66F5",
x"7EBB66B0",
x"7EE06663",
x"7EC26610",
x"7E7065B8",
x"7DFA6560",
x"7D76650E",
x"7CF764C9",
x"7C91649A",
x"7C506484",
x"7C3E6490",
x"7C5964BF",
x"7CA16511",
x"7D0B6584",
x"7D8E660E",
x"7E1E66A7",
x"7EAE673F",
x"7F3267CB",
x"7FA26841",
x"7FF96899",
x"803268CC",
x"804B68DF",
x"804468D5",
x"801D68B4",
x"7FDB6886",
x"7F806854",
x"7F136823",
x"7E9867F7",
x"7E1A67D5",
x"7DA067BC",
x"7D3467AA",
x"7CE0679D",
x"7CAE6794",
x"7CA16791",
x"7CBE6799",
x"7D0167AB",
x"7D6867CE",
x"7DE56804",
x"7E6C684C",
x"7EF168A4",
x"7F666904",
x"7FBF6962",
x"7FF469B0",
x"800469E5",
x"7FED69F7",
x"7FBA69E5",
x"7F7069AD",
x"7F1B6956",
x"7EC968ED",
x"7E86687F",
x"7E566817",
x"7E4567C5",
x"7E53678C",
x"7E816770",
x"7ECC676D",
x"7F2C677C",
x"7F9B678D",
x"800A6799",
x"806F6791",
x"80BB6773",
x"80E3673C",
x"80DC66EF",
x"80A06694",
x"802A6635",
x"7F7F65DE",
x"7EA46594",
x"7DA86560",
x"7C9A6541",
x"7B8E6534",
x"7A976531",
x"79C56531",
x"7927652D",
x"78C2651E",
x"789B6503",
x"78B064DF",
x"78F564B7",
x"795D6494",
x"79DC6481",
x"7A5D6486",
x"7ACE64A5",
x"7B1864DE",
x"7B2A6527",
x"7AEC6573",
x"7A4F65AE",
x"794265C1",
x"77BB6594",
x"75B56515",
x"73386437",
x"705162F3",
x"6D1A6150",
x"69B75F5D",
x"66525D36",
x"631C5AFD",
x"604158D9",
x"5DEC56F0",
x"5C3D5564",
x"5B485453",
x"5B1153C9",
x"5B8D53CC",
x"5CA45450",
x"5E34553F",
x"6013567A",
x"621757E1",
x"641D5950",
x"66035AAB",
x"67B55BDD",
x"692A5CD9",
x"6A615D9F",
x"6B5E5E38",
x"6C335EB1",
x"6CE95F1B",
x"6D945F84",
x"6E3B5FFA",
x"6EE5607E",
x"6F946111",
x"704661AB",
x"70F3623E",
x"719362BB",
x"721E6317",
x"728D6346",
x"72DB6346",
x"73066315",
x"731162BC",
x"73026246",
x"72DE61C2",
x"72AE613F",
x"727D60CB",
x"724F606E",
x"722D6035",
x"7217601E",
x"72106029",
x"72186053",
x"722D6093",
x"724B60E0",
x"72736135",
x"72A66188",
x"72E261D8",
x"732E6221",
x"738E6266",
x"740C62AD",
x"74AB62FC",
x"756F635C",
x"765B63D3",
x"7769646A",
x"78916523",
x"79C965F7",
x"7B0366E3",
x"7C2E67D6",
x"7D4268C5",
x"7E37699C",
x"7F096A4B",
x"7FBC6AC8",
x"805D6B0D",
x"80F36B1C",
x"818B6AF9",
x"822F6AB5",
x"82DF6A5E",
x"83986A03",
x"845069B5",
x"84F7697F",
x"85796962",
x"85C8695F",
x"85DB6972",
x"85AE6990",
x"854C69B1",
x"84CB69D2",
x"844469ED",
x"83D86A06",
x"83A46A1E",
x"83BE6A3F",
x"84316A6B",
x"84FB6AA3",
x"860B6AE6",
x"87466B2D",
x"88886B6F",
x"89AF6BA0",
x"8A9A6BB5",
x"8B356BAB",
x"8B796B7F",
x"8B696B38",
x"8B186AE5",
x"8AA16A96",
x"8A1D6A5B",
x"89A86A44",
x"89556A5B",
x"89296AA1",
x"89276B11",
x"89416B9D",
x"89666C33",
x"89866CBD",
x"898E6D2B",
x"89796D75",
x"89426D94",
x"88F36D8D",
x"889A6D6C",
x"88496D3F",
x"88116D16",
x"87FE6D00",
x"881A6D06",
x"885F6D28",
x"88C66D63",
x"893F6DAD",
x"89B76DF9",
x"8A1A6E3A",
x"8A596E62",
x"8A666E6B",
x"8A3E6E4D",
x"89DC6E09",
x"89426DA1",
x"88766D19",
x"87766C75",
x"86426BB4",
x"84D96ADB",
x"833469E6",
x"815168D5",
x"7F2B67A8",
x"7CC86662",
x"7A316507",
x"777763A1",
x"74B5623E",
x"720760E7",
x"6F8D5FAE",
x"6D685E9B",
x"6BAB5DB8",
x"6A6C5D07",
x"69AE5C8B",
x"696F5C40",
x"69A35C25",
x"6A375C33",
x"6B175C6D",
x"6C2E5CD2",
x"6D6F5D64",
x"6ECE5E2C",
x"70485F2F",
x"71DF6070",
x"739A61F2",
x"758363AD",
x"77A1659B",
x"79FC67B0",
x"7C9569D6",
x"7F6D6BFF",
x"827D6E19",
x"85BB7012",
x"891771E1",
x"8C84737E",
x"8FF274EA",
x"934D7626",
x"968A7737",
x"99977827",
x"9C6C78FB",
x"9EFD79BC",
x"A1487A6F",
x"A34B7B1C",
x"A50D7BC4",
x"A6947C6E",
x"A7F17D1C",
x"A9357DD0",
x"AA6E7E8C",
x"ABAF7F53",
x"AD058026",
x"AE778102",
x"B00781E1",
x"B1AC82BF",
x"B35A838F",
x"B4FE8446",
x"B68584D9",
x"B7DB853B",
x"B8F28563",
x"B9C2854C",
x"BA4D84F8",
x"BA9C8471",
x"BAC383C6",
x"BAD7830A",
x"BAF18256",
x"BB2581C6",
x"BB848170",
x"BC128166",
x"BCC981B0",
x"BD98824F",
x"BE678332",
x"BF168443",
x"BF898566",
x"BFA2867A",
x"BF548763",
x"BE998808",
x"BD7E8863",
x"BC1E8876",
x"BA9F884D",
x"B92F880A",
x"B7FE87C9",
x"B73A87B2",
x"B70487E0",
x"B76B8869",
x"B8718950",
x"BA018A90",
x"BBF48C0A",
x"BE188D9D",
x"C0338F1B",
x"C209905B",
x"C36A9135",
x"C42F9191",
x"C4449166",
x"C3AD90BB",
x"C27E8FA8",
x"C0DD8E52",
x"BEFC8CE6",
x"BD128B94",
x"BB548A85",
x"B9ED89DA",
x"B8F889A4",
x"B87E89E3",
x"B8778A85",
x"B8C68B6D",
x"B9448C6F",
x"B9C48D5C",
x"BA198E09",
x"BA228E50",
x"B9C98E1D",
x"B9118D6A",
x"B80C8C48",
x"B6E08AD3",
x"B5C0893C",
x"B4E487B9",
x"B4828681",
x"B4C085C5",
x"B5B685A9",
x"B760863F",
x"B9A28781",
x"BC468959",
x"BF088B97",
x"C19B8E01",
x"C3AF9059",
x"C505925D",
x"C57193D8",
x"C4E194A1",
x"C35E94A4",
x"C11393E5",
x"BE379276",
x"BB13907E",
x"B7ED8E2C",
x"B4FE8BB4",
x"B26D893C",
x"B04086E9",
x"AE6484C9",
x"ACAC82DD",
x"AAD18114",
x"A88E7F50",
x"A5A17D72",
x"A1D97B5B",
x"9D2778F5",
x"979B763C",
x"916D7339",
x"8AF07008",
x"848B6CD2",
x"7EAC69C7",
x"79B56714",
x"75F764E8",
x"739E6359",
x"72B56277",
x"7321623C",
x"74AD6295",
x"770D6365",
x"79F36487",
x"7D1165DE",
x"802E674C",
x"831E68BF",
x"85D36A30",
x"884F6B99",
x"8AA86CFF",
x"8CF66E69",
x"8F556FDC",
x"91D87157",
x"948B72D5",
x"976C7452",
x"9A6A75C7",
x"9D73772A",
x"A06B7878",
x"A33879AF",
x"A5C37AD4",
x"A7FD7BEB",
x"A9DC7CFE",
x"AB5D7E0F",
x"AC857F22",
x"AD5A8033",
x"ADEA813C",
x"AE42822F",
x"AE6B8301",
x"AE7583A3",
x"AE718412",
x"AE6B844D",
x"AE77845A",
x"AEA68449",
x"AF08842C",
x"AFAE841B",
x"B0A2842B",
x"B1ED846A",
x"B38B84E3",
x"B5758598",
x"B79B8681",
x"B9E6878F",
x"BC3888AE",
x"BE7289C8",
x"C0788AC8",
x"C22D8B9F",
x"C37E8C43",
x"C4608CB2",
x"C4D18CF1",
x"C4DB8D0E",
x"C4918D15",
x"C4098D18",
x"C3648D28",
x"C2BF8D4F",
x"C2328D95",
x"C1D38DFD",
x"C1AD8E80",
x"C1C78F16",
x"C2188FB5",
x"C2969053",
x"C32F90E7",
x"C3D09169",
x"C46791D5",
x"C4E4922E",
x"C5409273",
x"C57792A8",
x"C58B92D3",
x"C58592F7",
x"C56F9316",
x"C5579331",
x"C547934B",
x"C54A9363",
x"C56A937F",
x"C5A993A0",
x"C60993CC",
x"C68C940A",
x"C72C945E",
x"C7E294C9",
x"C8A9954C",
x"C97795DF",
x"CA419679",
x"CAFB9709",
x"CB9C9782",
x"CC1897D2",
x"CC6797EE",
x"CC8597CB",
x"CC729769",
x"CC3696CF",
x"CBDB9607",
x"CB749525",
x"CB10943F",
x"CAC9936A",
x"CAB092BF",
x"CAD7924E",
x"CB4A9224",
x"CC0C9249",
x"CD1B92BB",
x"CE6A9373",
x"CFE59463",
x"D1729579",
x"D2F7969D",
x"D45197B7",
x"D56598B0",
x"D6199970",
x"D65A99E8",
x"D61B9A0C",
x"D55B99D5",
x"D426994A",
x"D28C9872",
x"D0A7975E",
x"CE929620",
x"CC6594C7",
x"CA309360",
x"C7F591F2",
x"C5A99077",
x"C32D8EDF",
x"C0518D13",
x"BCE38AF3",
x"B8A68860",
x"B3718542",
x"AD25818A",
x"A5C87D3A",
x"9D777867",
x"94797337",
x"8B2C6DE8",
x"820B68BA",
x"799363FA",
x"723B5FED",
x"6C695CCD",
x"68635AC0",
x"664759D9",
x"660C5A10",
x"67825B45",
x"6A5F5D48",
x"6E445FDF",
x"72CB62C8",
x"779365C4",
x"7C4E689D",
x"80BB6B28",
x"84B46D4B",
x"88286EFA",
x"8B177037",
x"8D8A710D",
x"8F947190",
x"914571DA",
x"92AC71FF",
x"93D7721A",
x"94C97239",
x"9588726B",
x"961472B9",
x"96707321",
x"969E73A5",
x"96A8743B",
x"969474DC",
x"966D757B",
x"963F760C",
x"96187685",
x"960376DE",
x"96087710",
x"962F771C",
x"967C7705",
x"96EC76D0",
x"97787689",
x"981B763A",
x"98C275EF",
x"995D75B3",
x"99DC7590",
x"9A2E758C",
x"9A4A75AC",
x"9A2E75F1",
x"99E17658",
x"997676E2",
x"99047788",
x"98A87847",
x"98837916",
x"98AE79F1",
x"993B7ACE",
x"9A317BA5",
x"9B877C6B",
x"9D287D16",
x"9EF47D9E",
x"A0C67DF8",
x"A2787E1E",
x"A3E77E0B",
x"A4FD7DC3",
x"A5A77D47",
x"A5E67CA5",
x"A5C27BE7",
x"A54C7B1F",
x"A4987A5E",
x"A3C279B7",
x"A2E1793A",
x"A21078F5",
x"A16378F4",
x"A0F07937",
x"A0CC79C4",
x"A10A7A95",
x"A1B57BA0",
x"A2D77CD9",
x"A4717E32",
x"A6757F99",
x"A8D08100",
x"AB5D8256",
x"ADF1838C",
x"B05D8499",
x"B2708576",
x"B3FE861C",
x"B4EB868F",
x"B52C86D2",
x"B4C286E7",
x"B3C786DA",
x"B26086B3",
x"B0B9867A",
x"AF028635",
x"AD6785EC",
x"AC0885A2",
x"AAF4855A",
x"AA2C8514",
x"A9A884CC",
x"A9508482",
x"A90B8433",
x"A8C083DD",
x"A8598380",
x"A7D0831C",
x"A72682B8",
x"A66B8257",
x"A5B88202",
x"A52881C0",
x"A4DA8198",
x"A4E6818E",
x"A55A81A3",
x"A63581D6",
x"A76A821C",
x"A8D9826B",
x"AA5982B5",
x"ABBC82EB",
x"ACD68302",
x"AD7D82F1",
x"AD9C82B8",
x"AD298259",
x"AC3281E0",
x"AACA8156",
x"A91880CA",
x"A7428046",
x"A5667FCA",
x"A3987F53",
x"A1D77ED1",
x"A0127E2A",
x"9E277D44",
x"9BE67C02",
x"99257A4B",
x"95C27815",
x"91AE7561",
x"8CF77241",
x"87C96EDB",
x"826C6B62",
x"7D3A680E",
x"78976521",
x"74E662D2",
x"7275614F",
x"717960B4",
x"72036108",
x"74036241",
x"7748643B",
x"7B8466C9",
x"806269B5",
x"85836CC4",
x"8A916FBD",
x"8F467275",
x"936D74C7",
x"96E976A3",
x"99AF7802",
x"9BC278EA",
x"9D337968",
x"9E187993",
x"9E857982",
x"9E92794A",
x"9E5078FC",
x"9DCF78AA",
x"9D1B785A",
x"9C407810",
x"9B4B77CE",
x"9A437790",
x"99357755",
x"98297718",
x"972976D8",
x"963F7695",
x"956E7651",
x"94C17610",
x"943875DA",
x"93DA75B3",
x"93A8759F",
x"93A475A3",
x"93CD75C0",
x"942175F4",
x"949A763A",
x"952B768D",
x"95CB76E2",
x"96677731",
x"96F1776E",
x"975A7790",
x"97957793",
x"979A7772",
x"9763772C",
x"96F476C4",
x"9656763E",
x"959775A5",
x"94C574FE",
x"93F67454",
x"933973B1",
x"92A1731F",
x"923B72A6",
x"92117250",
x"92257220",
x"927A721D",
x"93077247",
x"93C3729D",
x"949C7319",
x"958073B0",
x"96597457",
x"971074FC",
x"978D7590",
x"97BE7601",
x"97957641",
x"970A7647",
x"961E760D",
x"94DC7597",
x"935674EF",
x"91A47423",
x"8FE47344",
x"8E397265",
x"8CBF719C",
x"8B9170F6",
x"8AC27083",
x"8A5F704B",
x"8A677051",
x"8AD67094",
x"8B9B7112",
x"8CA271C0",
x"8DD57295",
x"8F157385",
x"904F7485",
x"916D7583",
x"925F7674",
x"93177744",
x"939477EA",
x"93D57853",
x"93DD7879",
x"93B87857",
x"937177EC",
x"931B7743",
x"92C57668",
x"92837571",
x"92647478",
x"927B739A",
x"92D572F2",
x"937B729A",
x"947372A6",
x"95BB731C",
x"974973FC",
x"9912753B",
x"9AFE76C4",
x"9CF67875",
x"9EDA7A2D",
x"A0917BC4",
x"A1FD7D18",
x"A30C7E0B",
x"A3B37E88",
x"A3EE7E8A",
x"A3C57E12",
x"A3467D30",
x"A2877BFE",
x"A19E7A98",
x"A09F791D",
x"9F9277A6",
x"9E7B7647",
x"9D4B7508",
x"9BE673E5",
x"9A2C72D1",
x"97F671B3",
x"95187073",
x"917A6EF6",
x"8D0E6D26",
x"87DB6AF7",
x"81FE686C",
x"7BB26591",
x"753E6284",
x"6EF75F69",
x"693A5C6C",
x"645959BB",
x"609F577F",
x"5E3555DA",
x"5D3654E3",
x"5D96549E",
x"5F305505",
x"61CB5604",
x"651E577E",
x"68DB594D",
x"6CB15B4D",
x"705F5D5A",
x"73B45F58",
x"7690612E",
x"78EB62D2",
x"7ACC643F",
x"7C4E657C",
x"7D906690",
x"7EB8678A",
x"7FE96877",
x"813E6961",
x"82C96A4E",
x"848E6B41",
x"868A6C37",
x"88AD6D28",
x"8ADF6E0A",
x"8D076ED4",
x"8F106F76",
x"90DF6FEE",
x"92677035",
x"939B704D",
x"94777039",
x"94FD7005",
x"952E6FBD",
x"95126F6E",
x"94B46F26",
x"941B6EF0",
x"93526ED7",
x"92626ED8",
x"91566EF3",
x"903E6F26",
x"8F226F61",
x"8E156F9D",
x"8D256FCE",
x"8C5D6FEC",
x"8BCC6FF0",
x"8B766FD9",
x"8B5D6FAD",
x"8B806F6E",
x"8BD56F27",
x"8C4C6EE1",
x"8CD96EA1",
x"8D676E73",
x"8DE76E57",
x"8E4D6E4F",
x"8E8E6E5B",
x"8EAA6E79",
x"8EA16EA4",
x"8E7A6EDC",
x"8E3F6F1D",
x"8DFD6F64",
x"8DC26FAD",
x"8D976FF5",
x"8D87703A",
x"8D957073",
x"8DC3709D",
x"8E0B70B3",
x"8E6970AD",
x"8ECC708A",
x"8F2C704B",
x"8F796FF5",
x"8FA76F8F",
x"8FAC6F21",
x"8F836EBA",
x"8F2B6E62",
x"8EA56E21",
x"8DF96DFC",
x"8D316DF0",
x"8C566DF9",
x"8B736E09",
x"8A916E13",
x"89B76E0A",
x"88E36DE1",
x"88186D8F",
x"87536D12",
x"868D6C6B",
x"85C26BA1",
x"84EF6AC1",
x"841369D8",
x"832E68F2",
x"8243681B",
x"8159675B",
x"807766B4",
x"7FA16627",
x"7EE065B1",
x"7E38654C",
x"7DAD64F2",
x"7D4464A0",
x"7CFC6455",
x"7CDA6413",
x"7CDE63E0",
x"7D0463C6",
x"7D4E63CE",
x"7DB563FD",
x"7E32645A",
x"7EBB64E3",
x"7F446593",
x"7FBE665C",
x"801D672E",
x"805267F5",
x"8053689B",
x"801A690E",
x"7FA5693F",
x"7EF76926",
x"7E1768BC",
x"7D0A680A",
x"7BDC6717",
x"7A9365EF",
x"793164A1",
x"77B7633E",
x"762161CF",
x"746C6062",
x"728D5EFA",
x"70835D9B",
x"6E4A5C48",
x"6BE85B01",
x"696959C6",
x"66E2589C",
x"646C5788",
x"62275691",
x"603455C0",
x"5EB35525",
x"5DC054C7",
x"5D6F54B5",
x"5DCB54F3",
x"5ED25585",
x"60795669",
x"62A85797",
x"65445901",
x"68245A95",
x"6B275C3D",
x"6E245DE4",
x"70FC5F72",
x"739760D3",
x"75E561FD",
x"77DD62E8",
x"79876395",
x"7AEA640B",
x"7C1B6459",
x"7D2B6490",
x"7E3064C1",
x"7F3A64FF",
x"80526553",
x"817E65C8",
x"82BC665C",
x"8400670A",
x"853C67C5",
x"86606880",
x"875B6927",
x"882069B0",
x"88A76A0F",
x"88ED6A3D",
x"88F66A3E",
x"88CB6A17",
x"887969D5",
x"88116984",
x"87A06937",
x"873168F6",
x"86CD68CF",
x"867768C5",
x"862B68D6",
x"85E368FF",
x"85976935",
x"853C696F",
x"84CB69A3",
x"843C69C7",
x"839469D6",
x"82D369D4",
x"820A69C2",
x"814369AA",
x"80946994",
x"800D698A",
x"7FBF6997",
x"7FB869BB",
x"7FF969FA",
x"80836A4E",
x"81496AAD",
x"823B6B0F",
x"83416B65",
x"84426BA3",
x"85286BBF",
x"85DB6BB5",
x"864E6B83",
x"867A6B2B",
x"86606AB8",
x"860B6A35",
x"858969AE",
x"84EC6932",
x"844668CF",
x"83AA688D",
x"83276876",
x"82C4688D",
x"828768D1",
x"8270693E",
x"827E69CB",
x"82AD6A72",
x"82F66B23",
x"83526BD5",
x"83BE6C7C",
x"84346D0F",
x"84AC6D86",
x"85256DDE",
x"85946E16",
x"85F36E30",
x"86386E2E",
x"865D6E16",
x"865F6DEE",
x"86386DBA",
x"85EC6D7F",
x"85806D41",
x"85006D03",
x"84766CC8",
x"83F46C92",
x"83876C63",
x"833C6C41",
x"831F6C30",
x"83346C33",
x"83796C4E",
x"83EA6C80",
x"847D6CC8",
x"85206D20",
x"85C46D7D",
x"86536DD5",
x"86BC6E17",
x"86EF6E34",
x"86DC6E21",
x"867D6DD4",
x"85CE6D48",
x"84D36C82",
x"83976B89",
x"822A6A6D",
x"80A16942",
x"7F116819",
x"7D946703",
x"7C3B660E",
x"7B136544",
x"7A2364A3",
x"79666424",
x"78D363BE",
x"7855635F",
x"77D362F7",
x"77346277",
x"766361D3",
x"754C6106",
x"73EC6011",
x"72425EFD",
x"705F5DD7",
x"6E5C5CB5",
x"6C5B5BA6",
x"6A7F5AC2",
x"68EB5A17",
x"67BE59AE",
x"6711598C",
x"66EF59B3",
x"67585A1C",
x"68425ABD",
x"699E5B8A",
x"6B535C77",
x"6D455D78",
x"6F5E5E87",
x"71835F9B",
x"73A760B1",
x"75BE61C5",
x"77C562D6",
x"79BB63E6",
x"7BA364F2",
x"7D8365F9",
x"7F6266F7",
x"814167EC",
x"832368D5",
x"850769B2",
x"86ED6A83",
x"88CC6B48",
x"8A9F6C03",
x"8C606CB7",
x"8E036D65",
x"8F806E0D",
x"90CF6EAB",
x"91E96F40",
x"92C96FC5",
x"93717037",
x"93E37092",
x"942670D8",
x"94467108",
x"944D7127",
x"94497139",
x"943F7143",
x"94317144",
x"9412713A",
x"93D5711D",
x"935C70DF",
x"9288706F",
x"913B6FBD",
x"8F596EBA",
x"8CD86D61",
x"89B86BB2",
x"860E69C1",
x"820467A7",
x"7DD36587",
x"79BA6390",
x"75FC61E6",
x"72D660AF",
x"70766004",
x"6EF25FEA",
x"6E4B605C",
x"6E6D613F",
x"6F32626F",
x"706663C2",
x"71D2650B",
x"73426625",
x"748C66F3",
x"75936762",
x"764A6773",
x"76B1672E",
x"76D866A8",
x"76CF65FC",
x"76B06542",
x"768F6494",
x"767C6407",
x"768063A8",
x"769D637A",
x"76CB637C",
x"76FA63A3",
x"771A63E0",
x"77146423",
x"76D26459",
x"76426472",
x"755B645D",
x"741B6415",
x"72906398",
x"70D562ED",
x"6F116224",
x"6D796152",
x"6C456095",
x"6BB0600B",
x"6BEB5FD2",
x"6D196000",
x"6F4860A5",
x"726F61C5",
x"76696355",
x"7AFD653F",
x"7FE26760",
x"84C46994",
x"89536BB0",
x"8D4D6D8D",
x"907D6F0F",
x"92CA7023",
x"943470C1",
x"94CD70F2",
x"94C170C4",
x"943F7052",
x"937B6FB5",
x"92A76F0C",
x"91E46E68",
x"914E6DDB",
x"90E66D6B",
x"90AB6D17",
x"90886CD9",
x"906C6CA8",
x"903C6C7A",
x"8FEA6C48",
x"8F6D6C0D",
x"8EC36BCE",
x"8DF76B92",
x"8D1B6B5F",
x"8C436B44",
x"8B856B48",
x"8AF46B6F",
x"8A946BB4",
x"8A606C0A",
x"8A456C61",
x"8A226C9A",
x"89CB6C9D",
x"890D6C4B",
x"87B96B8D",
x"85A56A56",
x"82B868A1",
x"7EEB6677",
x"7A4E63EF",
x"75096127",
x"6F5C5E46",
x"69915B78",
x"63FD58E9",
x"5EF556BD",
x"5ABE5512",
x"579353FB",
x"5593537E",
x"54C75398",
x"551F5438",
x"56765544",
x"589956A4",
x"5B4A5835",
x"5E4A59D7",
x"61645B70",
x"64655CE9",
x"672A5E33",
x"69A05F45",
x"6BBD601B",
x"6D7F60B9",
x"6EF26129",
x"70206177",
x"711661AD",
x"71E161D6",
x"728961FC",
x"73146227",
x"73896258",
x"73E66290",
x"742F62C8",
x"746562FC",
x"7489631F",
x"749D632D",
x"74A46318",
x"74A162DC",
x"74976273",
x"748761DC",
x"7472611D",
x"74566039",
x"74345F3F",
x"74065E3B",
x"73C95D41",
x"737D5C60",
x"731E5BAB",
x"72B15B33",
x"72385B02",
x"71BA5B21",
x"713E5B8D",
x"70CE5C42",
x"706F5D32",
x"702B5E4B",
x"70055F76",
x"6FFC609D",
x"701461A9",
x"70486289",
x"7096632D",
x"70F66390",
x"716563B2",
x"71DD639B",
x"725B6355",
x"72D862ED",
x"73516276",
x"73C161F9",
x"74236186",
x"74746121",
x"74B160D0",
x"74D66095",
x"74E5606E",
x"74DF6058",
x"74C9604F",
x"74AB6050",
x"748D605C",
x"7476606E",
x"7470608A",
x"748260AE",
x"74AB60DC",
x"74F06114",
x"754E6158",
x"75BE61A7",
x"763A6201",
x"76BA6264",
x"773762CF",
x"77A7633E",
x"780663AA",
x"784B6411",
x"7875646F",
x"787D64BB",
x"786764F6",
x"7832651A",
x"77E5652A",
x"77866527",
x"771E6517",
x"76BE6501",
x"767364F0",
x"764A64ED",
x"764F64FF",
x"768F652A",
x"770B6573",
x"77C265D9",
x"78AD6655",
x"79BF66E0",
x"7AE56772",
x"7C0D67FD",
x"7D216877",
x"7E0E68DB",
x"7EC5691D",
x"7F3C693C",
x"7F6D6935",
x"7F586909",
x"7EFF68BA",
x"7E6D684C",
x"7DAF67C6",
x"7CD46730",
x"7BE86691",
x"7AFE65F6",
x"7A276566",
x"796D64EF",
x"78DD6498",
x"787C646C",
x"7845646C",
x"7834649B",
x"783764F3",
x"78386568",
x"782165E6",
x"77D8665C",
x"774466B0",
x"765566C8",
x"75046694",
x"73556603",
x"71566511",
x"6F2763C4",
x"6CE96229",
x"6ACB605D",
x"68F65E81",
x"67965CBB",
x"66C85B2F",
x"66A15A02",
x"6725594C",
x"684F591E",
x"6A05597A",
x"6C265A56",
x"6E8D5B9E",
x"71105D33",
x"73865EF7",
x"75D160C6",
x"77D36281",
x"79836410",
x"7ADB6562",
x"7BDE6670",
x"7C97673C",
x"7D1967CF",
x"7D726834",
x"7DB56877",
x"7DEF68A7",
x"7E2A68CE",
x"7E7068F0",
x"7EC46916",
x"7F25693B",
x"7F976962",
x"80176989",
x"80A469AB",
x"813F69C9",
x"81E869E5",
x"829A69FC",
x"83556A11",
x"84156A26",
x"84D66A3B",
x"85906A4F",
x"86386A62",
x"86C96A70",
x"87396A77",
x"87816A79",
x"879E6A70",
x"878E6A62",
x"87556A4F",
x"86F96A3E",
x"86866A35",
x"86076A3A",
x"858E6A51",
x"852A6A82",
x"84E56ACB",
x"84C96B2B",
x"84E26BA0",
x"852C6C20",
x"85AA6CA4",
x"86556D21",
x"87256D8F",
x"88106DE6",
x"890D6E23",
x"8A136E44",
x"8B186E4E",
x"8C176E48",
x"8D086E3B",
x"8DE56E31",
x"8EA76E37",
x"8F456E54",
x"8FB96E8D",
x"8FFA6EE5",
x"90006F57",
x"8FC66FDC",
x"8F4B7066",
x"8E9070E8",
x"8D9C714F",
x"8C80718C",
x"8B467192",
x"8A077157",
x"88D070D8",
x"87B87017",
x"86CB6F1E",
x"86136DFD",
x"85916CC7",
x"85466B93",
x"852C6A77",
x"853A6989",
x"856068D6",
x"8598686C",
x"85D66849",
x"86116868",
x"864568BC",
x"866D6934",
x"868B69BB",
x"86A46A3E",
x"86BB6AAD",
x"86DB6AFD",
x"870B6B30",
x"87566B44",
x"87C66B45",
x"88626B44",
x"892B6B4C",
x"8A226B6D",
x"8B3E6BB1",
x"8C746C1C",
x"8DB66CAE",
x"8EF36D62",
x"901A6E2E",
x"911A6F06",
x"91E96FDC",
x"928070A6",
x"92DF7157",
x"930471E8",
x"92F47252",
x"92B67292",
x"924E72A3",
x"91BE7286",
x"9108723A",
x"903171C4",
x"8F357127",
x"8E177069",
x"8CDA6F93",
x"8B7F6EAB",
x"8A076DB7",
x"88736CB8",
x"86BF6BB1",
x"84E56A9C",
x"82D8696D",
x"808C681E",
x"7DF366A4",
x"7B0764F9",
x"77C8631A",
x"74416111",
x"708A5EF0",
x"6CCE5CD0",
x"693E5AD3",
x"6614591A",
x"638757C6",
x"61CA56F5",
x"60FC56B8",
x"612D5712",
x"625157FE",
x"644D5964",
x"66EF5B29",
x"69FD5D29",
x"6D3A5F3F",
x"706C6149",
x"7365632B",
x"760464D3",
x"783F6634",
x"7A16674B",
x"7B98681B",
x"7CDE68AE",
x"7E00690D",
x"7F186944",
x"803B695F",
x"81746969",
x"82C86969",
x"84356969",
x"85B66970",
x"87436984",
x"88D069AB",
x"8A5869E9",
x"8BD06A3F",
x"8D386AAE",
x"8E8D6B37",
x"8FCC6BD5",
x"90F76C84",
x"92136D42",
x"93216E0A",
x"94266ED8",
x"95286FAB",
x"962C7082",
x"9733715A",
x"98407230",
x"99527302",
x"9A5F73CB",
x"9B607483",
x"9C487526",
x"9D0B75AC",
x"9D9F7612",
x"9E007654",
x"9E2B7678",
x"9E2C7683",
x"9E157685",
x"9E00768B",
x"9E0876A7",
x"9E4D76EC",
x"9EE97767",
x"9FE7781D",
x"A14F7912",
x"A3147A3A",
x"A5197B86",
x"A73C7CE3",
x"A9507E2F",
x"AB257F53",
x"AC958037",
x"AD8280C9",
x"ADE18100",
x"ADB580DB",
x"AD15806D",
x"AC267FC6",
x"AB147F02",
x"AA0E7E40",
x"A93C7D98",
x"A8BD7D1E",
x"A8A17CDD",
x"A8DF7CD7",
x"A9617CFF",
x"AA077D44",
x"AAA17D8C",
x"AB047DC0",
x"AB0A7DC9",
x"AA947D99",
x"A99A7D2C",
x"A81C7C86",
x"A62F7BB7",
x"A3F37AD4",
x"A18B79F1",
x"9F1F7926",
x"9CD67881",
x"9AC87809",
x"990B77BE",
x"97A97799",
x"96A2778B",
x"95F07783",
x"95887775",
x"95627755",
x"956E7720",
x"95A976D8",
x"96067685",
x"967D7631",
x"970475E8",
x"979275B0",
x"981D758C",
x"9894757B",
x"98EC7572",
x"99157567",
x"9908754A",
x"98BF7510",
x"983574B4",
x"97707433",
x"96787395",
x"955772E4",
x"941B7236",
x"92D27199",
x"91887121",
x"904D70DC",
x"8F2B70CD",
x"8E2B70EF",
x"8D577139",
x"8CB57197",
x"8C4671F4",
x"8C077234",
x"8BF17241",
x"8BF37209",
x"8BF7717C",
x"8BDD7094",
x"8B876F54",
x"8AD26DBF",
x"899F6BE6",
x"87DC69D9",
x"857F67AE",
x"8290657A",
x"7F2C6355",
x"7B7C6155",
x"77B85F8B",
x"741E5E0E",
x"70EF5CEC",
x"6E635C2F",
x"6CAA5BE3",
x"6BE25C0A",
x"6C145CA2",
x"6D3B5DA4",
x"6F3C5F04",
x"71F960B2",
x"7545629B",
x"78F964AB",
x"7CED66CE",
x"810768F2",
x"852E6B07",
x"89566D08",
x"8D796EEC",
x"919070B4",
x"95977265",
x"998A7400",
x"9D59758C",
x"A0F4770B",
x"A445787E",
x"A73079DE",
x"A99F7B23",
x"AB7B7C43",
x"ACB97D2F",
x"AD527DDA",
x"AD4F7E3C",
x"ACC67E51",
x"ABCF7E19",
x"AA917D9E",
x"A9327CED",
x"A7DA7C1C",
x"A6AE7B43",
x"A5C97A78",
x"A53D79D3",
x"A5157964",
x"A5507939",
x"A5E67956",
x"A6C879BD",
x"A7EA7A6A",
x"A93F7B56",
x"AABF7C75",
x"AC667DC1",
x"AE327F30",
x"B02C80BA",
x"B257825A",
x"B4B38405",
x"B73A85B5",
x"B9E38760",
x"BC9288F9",
x"BF2D8A71",
x"C18C8BC0",
x"C38C8CD8",
x"C5088DAF",
x"C5E58E43",
x"C6188E94",
x"C5A08EA7",
x"C4918E84",
x"C30B8E3C",
x"C13D8DDC",
x"BF5D8D73",
x"BD9F8D10",
x"BC368CBB",
x"BB468C7B",
x"BAEA8C55",
x"BB298C49",
x"BBFB8C55",
x"BD4C8C77",
x"BEFA8CAE",
x"C0DB8CF6",
x"C2CC8D4B",
x"C4A58DAB",
x"C6468E0E",
x"C7998E71",
x"C8928EC9",
x"C92F8F10",
x"C9728F38",
x"C9688F3C",
x"C9208F14",
x"C8A78EBE",
x"C80C8E39",
x"C75D8D8E",
x"C6A08CC5",
x"C5E08BEC",
x"C51F8B14",
x"C4608A4C",
x"C3A689A4",
x"C2F28925",
x"C24988D6",
x"C1AF88BB",
x"C12888CF",
x"C0BC890E",
x"C0708970",
x"C04A89E9",
x"C0508A74",
x"C0828B07",
x"C0E18B9D",
x"C1678C32",
x"C20B8CC5",
x"C2C28D52",
x"C3798DD6",
x"C41F8E4C",
x"C49E8EAA",
x"C4DB8EE5",
x"C4C48EF0",
x"C4448EBE",
x"C3508E43",
x"C1DE8D7A",
x"BFF48C5F",
x"BD9C8AFA",
x"BAEE8959",
x"B807878F",
x"B50B85B8",
x"B21983ED",
x"AF548245",
x"ACCD80CF",
x"AA8B7F94",
x"A8817E8A",
x"A6947D9E",
x"A4977CB3",
x"A2557BA0",
x"9F957A43",
x"9C247875",
x"97DC761F",
x"92AC7336",
x"8CA16FC5",
x"85E36BE9",
x"7EB567D1",
x"777263B4",
x"707C5FD5",
x"6A3B5C71",
x"650D59C3",
x"613857F0",
x"5EE9570B",
x"5E2A5712",
x"5EE557EB",
x"60E55970",
x"63DF5B6A",
x"677C5D9E",
x"6B5F5FD3",
x"6F3461DC",
x"72B46393",
x"75AD64E2",
x"780365C5",
x"79B26648",
x"7AC9667A",
x"7B636677",
x"7BAA665C",
x"7BC46641",
x"7BD8663B",
x"7C076655",
x"7C656694",
x"7CFD66F6",
x"7DCE6770",
x"7ECB67F9",
x"7FE26881",
x"80FA68FF",
x"81FC6965",
x"82D069AE",
x"836669D9",
x"83B469E8",
x"83B569E1",
x"837469C9",
x"82FD69AD",
x"82656991",
x"81C26980",
x"812F697C",
x"80C2698A",
x"808D69AA",
x"809B69D9",
x"80F36A14",
x"818E6A59",
x"82656AA1",
x"83656AE9",
x"84776B30",
x"85876B72",
x"867E6BB1",
x"874D6BEF",
x"87E76C2D",
x"884B6C6D",
x"88796CB1",
x"887A6CF9",
x"88606D3F",
x"883B6D83",
x"881B6DBE",
x"88116DEC",
x"88276E09",
x"88626E16",
x"88C26E12",
x"89416E05",
x"89D66DF3",
x"8A796DEB",
x"8B1B6DF5",
x"8BB66E1C",
x"8C426E62",
x"8CB96ECD",
x"8D1D6F57",
x"8D6A6FF8",
x"8DA870A4",
x"8DD9714D",
x"8E0171E4",
x"8E27725C",
x"8E4972AF",
x"8E7072D5",
x"8E9A72D0",
x"8EC872A1",
x"8EF97255",
x"8F2971EF",
x"8F52717C",
x"8F6D7100",
x"8F737085",
x"8F5C700A",
x"8F216F96",
x"8EC16F29",
x"8E3E6EC5",
x"8D9E6E6E",
x"8CED6E23",
x"8C396DE8",
x"8B936DBF",
x"8B066DA9",
x"8A9E6DA1",
x"8A626DA7",
x"8A506DB3",
x"8A646DBB",
x"8A976DBD",
x"8AD96DAE",
x"8B246D8F",
x"8B696D5C",
x"8BA46D1C",
x"8BD26CD2",
x"8BF36C89",
x"8C096C47",
x"8C176C14",
x"8C226BF5",
x"8C286BE8",
x"8C286BEC",
x"8C206BF9",
x"8C076C09",
x"8BDC6C10",
x"8B9A6C0A",
x"8B446BF3",
x"8ADA6BCA",
x"8A646B93",
x"89E96B55",
x"896F6B14",
x"88F76AD7",
x"887E6A9E",
x"87FC6A66",
x"875B6A28",
x"868369D4",
x"8558695B",
x"83BB68AA",
x"819667B1",
x"7ED36668",
x"7B7464CB",
x"778362E3",
x"731E60C3",
x"6E735E84",
x"69BC5C48",
x"653D5A32",
x"61355866",
x"5DE65701",
x"5B7F5619",
x"5A2355B8",
x"59DE55DD",
x"5AA6567D",
x"5C5E5782",
x"5ED858D0",
x"61DF5A47",
x"65345BCB",
x"68A05D3F",
x"6BEF5E8E",
x"6EFA5FAE",
x"71AD609A",
x"73F96155",
x"75E561E9",
x"777D6268",
x"78D662E0",
x"7A076365",
x"7B2A6403",
x"7C4E64C6",
x"7D8065B2",
x"7EC966C6",
x"802567FC",
x"818D6945",
x"82F46A94",
x"844E6BD8",
x"858A6D00",
x"86A06E00",
x"87846ECD",
x"88386F64",
x"88BE6FC4",
x"891F6FF3",
x"896C6FFA",
x"89AE6FE2",
x"89F76FB7",
x"8A4F6F80",
x"8ABE6F48",
x"8B406F13",
x"8BD06EE4",
x"8C636EBD",
x"8CEA6EA1",
x"8D596E92",
x"8DA56E96",
x"8DCB6EB1",
x"8DCF6EEE",
x"8DBE6F51",
x"8DA86FE2",
x"8DA570A1",
x"8DCC718D",
x"8E32729C",
x"8EE673BE",
x"8FEE74E1",
x"914C75F1",
x"92F376DA",
x"94D2778D",
x"96D27801",
x"98DC7832",
x"9AD67826",
x"9CA877EA",
x"9E3D778D",
x"9F8A7723",
x"A07D76B7",
x"A115765A",
x"A14D760D",
x"A12B75D7",
x"A0B675B0",
x"9FFD7593",
x"9F127578",
x"9E0D7557",
x"9D04752F",
x"9C1174FB",
x"9B4C74BE",
x"9AC67480",
x"9A8B7446",
x"9A9F7416",
x"9AFE73F8",
x"9B9A73EF",
x"9C6073FE",
x"9D397423",
x"9E0D745E",
x"9EC674AC",
x"9F527506",
x"9FA4756B",
x"9FB975D5",
x"9F957640",
x"9F3F76A7",
x"9EC37705",
x"9E2E7755",
x"9D8B7790",
x"9CE777B2",
x"9C4677B3",
x"9BA8778C",
x"9B0D773A",
x"9A6F76BD",
x"99C57612",
x"990B7541",
x"98427451",
x"9767734D",
x"96867248",
x"95A57152",
x"94D77080",
x"942B6FE4",
x"93AB6F8A",
x"93626F7F",
x"93506FC0",
x"93707044",
x"93B670FE",
x"940E71D2",
x"946072A7",
x"949A7361",
x"94A573E5",
x"94777421",
x"940B740D",
x"936373A9",
x"928772FF",
x"91807220",
x"9058711F",
x"8F157012",
x"8DB86F05",
x"8C396E02",
x"8A8B6D0A",
x"88A46C14",
x"86716B13",
x"83EF69FA",
x"811E68BB",
x"7E0D6751",
x"7AD865BC",
x"77A36407",
x"749E6248",
x"71FA609A",
x"6FE65F1A",
x"6E865DE6",
x"6DF55D1A",
x"6E375CC8",
x"6F475CF6",
x"710C5DA4",
x"73605EC6",
x"761B6046",
x"790E620D",
x"7C1063FA",
x"7EFA65F5",
x"81B267DF",
x"842B69A6",
x"86606B3A",
x"88536C93",
x"8A136DAD",
x"8BAC6E8F",
x"8D2E6F3E",
x"8EA76FC7",
x"901B7034",
x"91937092",
x"930570E9",
x"946F7141",
x"95C2719D",
x"96F671FF",
x"98007265",
x"98D972CD",
x"99807334",
x"99FA739A",
x"9A4F7400",
x"9A907467",
x"9AC974D2",
x"9B10754B",
x"9B7075D2",
x"9BF6766F",
x"9CA97723",
x"9D8A77EB",
x"9E9578C3",
x"9FC279A5",
x"A10A7A8B",
x"A2637B6E",
x"A3C57C49",
x"A52C7D19",
x"A6977DE0",
x"A8087EA2",
x"A9827F60",
x"AB0A8020",
x"AC9C80E4",
x"AE3A81AB",
x"AFDF826E",
x"B17D8329",
x"B30783D2",
x"B46E8460",
x"B5A284CD",
x"B6958517",
x"B73F853B",
x"B79C853F",
x"B7B5852B",
x"B795850A",
x"B74F84E7",
x"B6FB84D0",
x"B6B384CC",
x"B69284E3",
x"B6AC8518",
x"B70F856E",
x"B7C385E3",
x"B8C68673",
x"BA0E8719",
x"BB8987D2",
x"BD298895",
x"BED78962",
x"C0848A2F",
x"C2268AFD",
x"C3B68BC8",
x"C5378C90",
x"C6B08D53",
x"C8278E16",
x"C9A38ED6",
x"CB238F98",
x"CCA39059",
x"CE129114",
x"CF5A91C2",
x"D05E9259",
x"D0FF92CB",
x"D1239304",
x"D0B492F9",
x"CFAA929A",
x"CE0891E0",
x"CBDD90CC",
x"C9478F67",
x"C6678DC5",
x"C3678BFD",
x"C06B8A31",
x"BD968883",
x"BB058714",
x"B8C98600",
x"B6EE8559",
x"B57B852C",
x"B4718576",
x"B3CE8629",
x"B38E872F",
x"B3A6886C",
x"B40B89BB",
x"B4A98AF9",
x"B56A8C07",
x"B62F8CC9",
x"B6D98D2B",
x"B7498D24",
x"B7678CB6",
x"B7208BEF",
x"B6748AE3",
x"B57089B1",
x"B42F8876",
x"B2D78753",
x"B18E8663",
x"B07785B6",
x"AFA68552",
x"AF1B8528",
x"AEBD8522",
x"AE5A8518",
x"ADB084DD",
x"AC748440",
x"AA5C8319",
x"A72C8146",
x"A2CD7EBD",
x"9D407B81",
x"96B677AF",
x"8F7C7375",
x"87FA6F12",
x"80AE6AC8",
x"7A0E66DC",
x"74836389",
x"705F60FA",
x"6DC95F49",
x"6CCB5E7D",
x"6D455E84",
x"6EFA5F41",
x"719E6088",
x"74DC622E",
x"78626401",
x"7BED65DF",
x"7F4F67A5",
x"826D6947",
x"853E6AB8",
x"87CC6C02",
x"8A2B6D2B",
x"8C706E44",
x"8EAE6F59",
x"90ED707A",
x"933471AB",
x"957472F1",
x"979F7446",
x"99A175A0",
x"9B6376F5",
x"9CD27839",
x"9DE3795B",
x"9E957A54",
x"9EF37B1B",
x"9F0E7BB0",
x"9F017C12",
x"9EED7C47",
x"9EF37C59",
x"9F2F7C4D",
x"9FB87C30",
x"A09E7C08",
x"A1DF7BE0",
x"A3737BBA",
x"A5437BA0",
x"A7337B93",
x"A91C7B98",
x"AADC7BB0",
x"AC4C7BE0",
x"AD527C26",
x"ADDE7C85",
x"ADED7CF8",
x"AD897D7E",
x"ACCD7E11",
x"ABD97EAC",
x"AAD97F49",
x"A9FB7FE6",
x"A96B8082",
x"A949811E",
x"A9A981BB",
x"AA8F825D",
x"ABF08308",
x"ADAC83BF",
x"AFA0847E",
x"B1A18540",
x"B3828601",
x"B52286B2",
x"B66A874A",
x"B75487BF",
x"B7EE880B",
x"B850882E",
x"B89E882F",
x"B8FF881B",
x"B9998803",
x"BA8887F9",
x"BBD98812",
x"BD88885C",
x"BF8688DD",
x"C1B38998",
x"C3E88A81",
x"C5FB8B88",
x"C7C98C97",
x"C9328D93",
x"CA298E66",
x"CAAC8EFD",
x"CAC78F4E",
x"CA938F55",
x"CA2C8F1D",
x"C9B38EB5",
x"C9448E35",
x"C8F48DB5",
x"C8CD8D4C",
x"C8D18D0E",
x"C8F78D03",
x"C9288D2E",
x"C94C8D83",
x"C9498DEF",
x"C9018E5D",
x"C8628EB1",
x"C7628ED6",
x"C5FB8EB8",
x"C4398E52",
x"C2308DA5",
x"BFFF8CBF",
x"BDC78BB6",
x"BBAF8AA5",
x"B9D689A8",
x"B85988D6",
x"B7468842",
x"B6A387F1",
x"B66487E0",
x"B6718801",
x"B6A8883F",
x"B6E48881",
x"B6FE88AE",
x"B6D388AE",
x"B64F8877",
x"B5648801",
x"B4188750",
x"B27A866E",
x"B0A1856A",
x"AEAB8452",
x"ACAF8331",
x"AABC820B",
x"A8D980E3",
x"A6F57FAF",
x"A4FD7E5E",
x"A2C77CE0",
x"A02F7B23",
x"9D10791B",
x"994D76C1",
x"94E3741F",
x"8FDD7140",
x"8A606E41",
x"84A76B45",
x"7EFA6872",
x"79AB65ED",
x"750663D9",
x"714F624E",
x"6EB76159",
x"6D5460FC",
x"6D236129",
x"6E0661C9",
x"6FCC62BC",
x"723763E0",
x"75006510",
x"77E56630",
x"7AAE672B",
x"7D3467F6",
x"7F636891",
x"8138690A",
x"82C26970",
x"841E69DC",
x"856D6A61",
x"86D16B13",
x"88636BFD",
x"8A356D20",
x"8C4C6E75",
x"8EA16FEF",
x"911E7176",
x"93AA72F8",
x"9627745E",
x"98797597",
x"9A8A769C",
x"9C4B776A",
x"9DB87806",
x"9ED7787E",
x"9FB278DB",
x"A05A7930",
x"A0E17988",
x"A15A79EA",
x"A1D27A57",
x"A2527AD0",
x"A2E67B4B",
x"A3917BC3",
x"A4577C2D",
x"A53F7C85",
x"A64C7CC7",
x"A7847CF5",
x"A8EA7D14",
x"AA847D2D",
x"AC507D4C",
x"AE4A7D7E",
x"B06E7DCD",
x"B2AD7E44",
x"B4FD7EE8",
x"B74F7FBC",
x"B99980C2",
x"BBD681F4",
x"BE01834D",
x"C01E84C3",
x"C22C864C",
x"C42D87DA",
x"C61F895F",
x"C7FA8ACA",
x"C9AD8C0D",
x"CB288D18",
x"CC4E8DDD",
x"CD0E8E53",
x"CD548E76",
x"CD188E43",
x"CC5E8DC5",
x"CB378D07",
x"C9C28C1A",
x"C81F8B13",
x"C6788A04",
x"C4F18904",
x"C3A58821",
x"C2A58763",
x"C1F186CD",
x"C17E865E",
x"C136860F",
x"C0FC85D4",
x"C0B685A2",
x"C04E856E",
x"BFB68535",
x"BEEE84F0",
x"BE0284A7",
x"BD04845C",
x"BC0F841C",
x"BB3C83F3",
x"BAA183EA",
x"BA44840A",
x"BA298454",
x"BA4084C5",
x"BA6E8550",
x"BA9385E6",
x"BA8C866E",
x"BA3686CF",
x"B97786F3",
x"B84586C3",
x"B6A08636",
x"B49F854A",
x"B263840B",
x"B01B828F",
x"ADFA80F7",
x"AC367F6B",
x"AAFA7E15",
x"AA647D16",
x"AA807C86",
x"AB437C75",
x"AC8E7CD9",
x"AE307D9E",
x"AFF07E9F",
x"B18F7FB0",
x"B2D480AC",
x"B3948168",
x"B3B681CD",
x"B33981D3",
x"B2338181",
x"B0C680ED",
x"AF228037",
x"AD777F82",
x"ABEA7EEE",
x"AA917E88",
x"A96E7E56",
x"A86D7E47",
x"A7677E41",
x"A62B7E1E",
x"A4877DB3",
x"A24D7CDE",
x"9F667B88",
x"9BC979A8",
x"978D7747",
x"92D97485",
x"8DE97188",
x"89046E80",
x"846F6B9E",
x"80676910",
x"7D2066F5",
x"7AB46560",
x"7931645A",
x"789063DC",
x"78BE63D5",
x"799B6432",
x"7B0764DC",
x"7CE065BB",
x"7F0666BC",
x"815C67D2",
x"83CE68F0",
x"86466A10",
x"88B96B2E",
x"8B1E6C4B",
x"8D6D6D65",
x"8FA76E7F",
x"91CE6F9C",
x"93E770C0",
x"95FD71EF",
x"981B732B",
x"9A4D747C",
x"9C9B75E1",
x"9F07775D",
x"A19178EB",
x"A42E7A8B",
x"A6D27C32",
x"A9677DD7",
x"ABDC7F6E",
x"AE1B80EB",
x"B0158242",
x"B1C08367",
x"B3178453",
x"B4178502",
x"B4C78573",
x"B52E85A8",
x"B55485A7",
x"B5448578",
x"B5088527",
x"B4A884BC",
x"B4308446",
x"B3B083CD",
x"B336835E",
x"B2D68300",
x"B2A182BB",
x"B2AB8291",
x"B3028287",
x"B3B2829B",
x"B4BA82CD",
x"B6188318",
x"B7B78377",
x"B98583E6",
x"BB64845A",
x"BD3584D3",
x"BED78546",
x"C03385B1",
x"C133860F",
x"C1CD865E",
x"C1FF869C",
x"C1CD86C6",
x"C14386DC",
x"C07586DA",
x"BF7786C0",
x"BE5E868E",
x"BD438643",
x"BC3885E0",
x"BB498568",
x"BA8284E4",
x"B9EB8456",
x"B98183CC",
x"B943834D",
x"B92882E6",
x"B92682A2",
x"B935828A",
x"B94A829F",
x"B95E82E7",
x"B970835C",
x"B97B83F6",
x"B98484A8",
x"B98B8566",
x"B9988621",
x"B9AD86CA",
x"B9CD8757",
x"B9F587C2",
x"BA228803",
x"BA4A881D",
x"BA638811",
x"BA5D87E2",
x"BA2C8794",
x"B9C3872B",
x"B91986A9",
x"B82B860E",
x"B6F88557",
x"B5898487",
x"B3ED839E",
x"B233829C",
x"B074818E",
x"AEC68078",
x"AD3D7F6B",
x"ABF37E77",
x"AAEE7DA5",
x"AA3B7D04",
x"A9D47C99",
x"A9B57C65",
x"A9C67C63",
x"A9F37C84",
x"AA1E7CB6",
x"AA2E7CE8",
x"AA077D06",
x"A99B7D05",
x"A8E17CDA",
x"A7DD7C85",
x"A6997C0F",
x"A5277B82",
x"A39B7AEE",
x"A20A7A60",
x"A07D79DE",
x"9EF4796B",
x"9D6478FB",
x"9BB3787C",
x"99BE77D5",
x"975D76EB",
x"946A759F",
x"90CE73DF",
x"8C7971A0",
x"877A6EE6",
x"81F36BC5",
x"7C1B685E",
x"763B64D8",
x"70A46164",
x"6BA65E35",
x"67855B71",
x"6473593C",
x"628C57A5",
x"61CC56B3",
x"621C5660",
x"63475697",
x"6512573D",
x"6738583A",
x"697F5971",
x"6BAD5AC9",
x"6DA35C31",
x"6F4B5D9A",
x"70A45EFD",
x"71BC6056",
x"72A861A5",
x"737D62E6",
x"74536417",
x"753C6535",
x"763E663B",
x"775C6723",
x"788E67E8",
x"79CC6884",
x"7B0A68FA",
x"7C3C6948",
x"7D5B6976",
x"7E62698A",
x"7F526990",
x"802D6991",
x"80F6699D",
x"81B169BA",
x"825F69ED",
x"82FE6A3E",
x"838B6AA8",
x"84006B26",
x"84586BAE",
x"848A6C37",
x"84956CB0",
x"847C6D0D",
x"84416D45",
x"83ED6D4E",
x"838E6D26",
x"83326CCF",
x"82EC6C4F",
x"82C86BB4",
x"82D26B0C",
x"83136A69",
x"838D69DE",
x"843F6977",
x"85216947",
x"862C6952",
x"8752699D",
x"88886A24",
x"89C16AE1",
x"8AF06BC5",
x"8C106CBE",
x"8D176DB8",
x"8E036EA0",
x"8ECD6F61",
x"8F796FEF",
x"90007041",
x"90667057",
x"90A87037",
x"90C56FF0",
x"90BE6F96",
x"90936F3D",
x"90436EF9",
x"8FD36EDC",
x"8F466EEF",
x"8E9F6F35",
x"8DE96FA6",
x"8D2A7034",
x"8C6C70CB",
x"8BBB7158",
x"8B2271C7",
x"8AAE7209",
x"8A66721C",
x"8A5271FE",
x"8A7471BA",
x"8ACE7164",
x"8B58710A",
x"8C0970C3",
x"8CD6709A",
x"8DAF709D",
x"8E8670C8",
x"8F497116",
x"8FEC717B",
x"906371E2",
x"90A8723A",
x"90B5726F",
x"908A7276",
x"90257244",
x"8F8D71D8",
x"8EC57139",
x"8DD3706F",
x"8CC16F88",
x"8B986E96",
x"8A696DAA",
x"893F6CD2",
x"882E6C1D",
x"87466B93",
x"86986B38",
x"862F6B0F",
x"86136B10",
x"86426B37",
x"86B86B79",
x"87656BC8",
x"88386C1A",
x"891B6C62",
x"89F96C9A",
x"8ABF6CBB",
x"8B606CC7",
x"8BD56CC2",
x"8C206CB4",
x"8C406CA7",
x"8C406CA3",
x"8C246CAB",
x"8BEA6CC2",
x"8B936CE1",
x"8B106CF9",
x"8A536CF9",
x"89486CCB",
x"87DB6C58",
x"85FD6B93",
x"83AA6A6F",
x"80E568F0",
x"7DC46723",
x"7A66651E",
x"76F66300",
x"73A760ED",
x"70AB5F08",
x"6E335D74",
x"6C625C48",
x"6B525B90",
x"6B095B50",
x"6B7C5B7E",
x"6C945C0A",
x"6E285CDC",
x"700F5DD7",
x"72175EE4",
x"74165FED",
x"75E860E2",
x"777361B5",
x"78B06268",
x"799D62FC",
x"7A4B6377",
x"7ACE63E6",
x"7B416455",
x"7BBE64CE",
x"7C5E655E",
x"7D2F660A",
x"7E3B66D6",
x"7F8067C1",
x"80F368C7",
x"828669DE",
x"84226AFC",
x"85B66C17",
x"872C6D24",
x"88796E1D",
x"89946EF9",
x"8A7D6FB5",
x"8B3B7055",
x"8BD670DA",
x"8C5F7145",
x"8CE0719D",
x"8D6971E5",
x"8E01721F",
x"8EAB724A",
x"8F647266",
x"902B7278",
x"90F4727C",
x"91B8727C",
x"9271727F",
x"931D728F",
x"93BE72BB",
x"945C7310",
x"9504739A",
x"95C8745F",
x"96B57560",
x"97D8768F",
x"993577E1",
x"9ACD793C",
x"9C957A84",
x"9E777B9F",
x"A0597C74",
x"A2217CF2",
x"A3AF7D12",
x"A4F17CD7",
x"A5D77C4D",
x"A6617B8B",
x"A6957AA9",
x"A68879C6",
x"A65378F8",
x"A6127856",
x"A5DD77E7",
x"A5C977B2",
x"A5DD77AD",
x"A61B77D0",
x"A6737809",
x"A6D27848",
x"A7227882",
x"A74C78A9",
x"A73E78BD",
x"A6F178C1",
x"A66A78BC",
x"A5B578B6",
x"A4E778BC",
x"A41E78D4",
x"A3737905",
x"A2FB794A",
x"A2C9799F",
x"A2DC79F8",
x"A32C7A49",
x"A3A97A7F",
x"A43B7A91",
x"A4C27A75",
x"A5257A26",
x"A54D79A8",
x"A52978FF",
x"A4B17837",
x"A3E4775D",
x"A2CC767E",
x"A17075A6",
x"9FE174DC",
x"9E2F7429",
x"9C69738B",
x"9A9E7302",
x"98DC728D",
x"97317229",
x"95A971D4",
x"9452718D",
x"9336715A",
x"925C713B",
x"91C37137",
x"9169714D",
x"9140717C",
x"913971C3",
x"913B7216",
x"9131726C",
x"910472B6",
x"90A872E8",
x"901772F9",
x"8F5672E1",
x"8E7672A1",
x"8D8D7240",
x"8CB471C7",
x"8C037143",
x"8B8970C3",
x"8B45704D",
x"8B2A6FE6",
x"8B1B6F8A",
x"8AF16F2D",
x"8A7D6EBE",
x"89936E26",
x"880D6D52",
x"85DB6C31",
x"82FC6ABB",
x"7F8468F2",
x"7BA066E2",
x"778464A3",
x"73756252",
x"6FB06011",
x"6C705E03",
x"69E15C43",
x"681B5AE9",
x"672959FD",
x"66FD5984",
x"67825975",
x"689359C3",
x"6A0C5A5D",
x"6BC25B32",
x"6D975C2E",
x"6F6D5D45",
x"71305E6D",
x"72D15F9D",
x"744F60D0",
x"75AE6203",
x"76F56331",
x"78306458",
x"796F6572",
x"7AC1667A",
x"7C37676C",
x"7DD66845",
x"7FA86903",
x"81A869AA",
x"83CC6A38",
x"86006AB7",
x"882B6B27",
x"8A346B90",
x"8BFE6BF5",
x"8D776C58",
x"8E906CBB",
x"8F436D1E",
x"8F9D6D7F",
x"8FAC6DDC",
x"8F8A6E33",
x"8F506E7F",
x"8F1A6EBE",
x"8EF66EEE",
x"8EF06F0A",
x"8F066F10",
x"8F2C6F00",
x"8F536ED8",
x"8F666E9A",
x"8F536E48",
x"8F116DE9",
x"8E9E6D83",
x"8E016D1E",
x"8D4C6CC4",
x"8C946C7A",
x"8BF36C4B",
x"8B796C34",
x"8B366C38",
x"8B2E6C54",
x"8B596C80",
x"8BA56CB4",
x"8BFD6CE8",
x"8C486D13",
x"8C6F6D31",
x"8C606D3E",
x"8C156D38",
x"8B936D24",
x"8AE06D08",
x"8A156CE5",
x"89466CC4",
x"888D6CAB",
x"87FD6CA0",
x"87A86CA4",
x"87966CBD",
x"87C66CE9",
x"88356D2A",
x"88D86D7C",
x"899F6DDC",
x"8A7C6E47",
x"8B5C6EB4",
x"8C316F1C",
x"8CEC6F76",
x"8D836FBB",
x"8DEA6FE4",
x"8E206FEB",
x"8E1B6FCE",
x"8DE26F92",
x"8D766F38",
x"8CE36ED1",
x"8C386E65",
x"8B876E05",
x"8AE26DBB",
x"8A596D93",
x"89FE6D92",
x"89D96DB7",
x"89E76DF9",
x"8A226E4F",
x"8A7A6EA9",
x"8AD86EF2",
x"8B246F1D",
x"8B466F1A",
x"8B2C6EE2",
x"8AC86E75",
x"8A186DD7",
x"89256D13",
x"87FD6C3D",
x"86B76B63",
x"856D6A9C",
x"843969F3",
x"83326976",
x"8265692B",
x"81DC690E",
x"8196691A",
x"818D6944",
x"81B1697F",
x"81F369BB",
x"823F69ED",
x"82846A0D",
x"82AF6A11",
x"82B569F9",
x"828D69C5",
x"82326976",
x"81A26910",
x"80E06894",
x"7FED6806",
x"7ED26763",
x"7D9166AE",
x"7C3265E2",
x"7ABD6500",
x"79346409",
x"77A06301",
x"760461ED",
x"746A60D8",
x"72D95FCB",
x"715B5ECF",
x"6FFC5DF1",
x"6ECC5D3C",
x"6DDB5CB3",
x"6D385C5D",
x"6CF55C39",
x"6D1E5C46",
x"6DBF5C84",
x"6EDB5CF1",
x"706F5D8D",
x"72765E59",
x"74E55F5A",
x"77AA6098",
x"7AB7621A",
x"7DFD63E5",
x"816F65FA",
x"85016859",
x"88B16AF7",
x"8C746DC5",
x"904970AD",
x"94267395",
x"98047661",
x"9BCF78F9",
x"9F737B46",
x"A2D77D3A",
x"A5E07ECF",
x"A8738002",
x"AA7A80E1",
x"ABE88178",
x"ACBC81D6",
x"ACFB820C",
x"ACB98226",
x"AC12822C",
x"AB258222",
x"AA148208",
x"A8F881D7",
x"A7EB818B",
x"A6FA811E",
x"A622808E",
x"A5607FDA",
x"A4A57F07",
x"A3E07E1C",
x"A3017D22",
x"A1FB7C22",
x"A0C97B25",
x"9F6E7A2F",
x"9DF77944",
x"9C777867",
x"9B047795",
x"99B876CB",
x"98AC760C",
x"97F17558",
x"979574B6",
x"979D742C",
x"980073C3",
x"98B27386",
x"99A2737E",
x"9AB673AA",
x"9BD5740D",
x"9CE474A0",
x"9DCD7554",
x"9E7B7619",
x"9EE276DD",
x"9EFB778C",
x"9EC97818",
x"9E547874",
x"9DAE789D",
x"9CEA7898",
x"9C227868",
x"9B70781D",
x"9AE777C4",
x"9A9C776A",
x"9A977718",
x"9AD776D5",
x"9B5976A9",
x"9C0B7690",
x"9CDA7689",
x"9DAF7696",
x"9E7A76B3",
x"9F2976E5",
x"9FB97731",
x"A02C779D",
x"A08B782D",
x"A0E678E5",
x"A14D79C4",
x"A1CF7AC0",
x"A2737BCA",
x"A3367CCE",
x"A40A7DB2",
x"A4D97E5D",
x"A5847EB9",
x"A5EE7EB7",
x"A5FE7E53",
x"A59F7D91",
x"A4CF7C81",
x"A3987B3D",
x"A21279E4",
x"A05F7895",
x"9EA5776B",
x"9D0A767E",
x"9BAC75D7",
x"9A9F7576",
x"99E77554",
x"9979755E",
x"993B757B",
x"990E7593",
x"98CD758F",
x"9858755B",
x"979274EE",
x"966E7443",
x"94EA735C",
x"93107245",
x"90F4710C",
x"8EB56FC1",
x"8C716E75",
x"8A436D34",
x"88436C0C",
x"867C6B03",
x"84EF6A1A",
x"8394694E",
x"82566896",
x"811A67E9",
x"7FBF6738",
x"7E256676",
x"7C346594",
x"79D6648A",
x"77046352",
x"73C561EC",
x"702A6059",
x"6C515EA9",
x"68605CE7",
x"64895B29",
x"60F25981",
x"5DC85801",
x"5B2A56BA",
x"592D55B9",
x"57DE5502",
x"573B5496",
x"5737546E",
x"57C45482",
x"58C854C6",
x"5A30552B",
x"5BE555A5",
x"5DD2562E",
x"5FE656BD",
x"62135751",
x"644857EA",
x"6676588B",
x"688D5938",
x"6A7D59F3",
x"6C355ABD",
x"6DA95B98",
x"6ECE5C7E",
x"6FA15D6C",
x"70285E59",
x"70705F3F",
x"70896018",
x"708960DD",
x"7086618D",
x"70936222",
x"70BB629F",
x"71046306",
x"716D6358",
x"71E96397",
x"726C63C6",
x"72E563E8",
x"734563FD",
x"7384640A",
x"73A1640D",
x"73A0640B",
x"73896407",
x"736D6403",
x"735C6404",
x"73666410",
x"73966425",
x"73F06446",
x"74766476",
x"752064B2",
x"75E264F7",
x"76B16546",
x"777D659A",
x"783C65F3",
x"78E5664E",
x"797266AA",
x"79E06703",
x"7A346759",
x"7A7067A5",
x"7A9E67E8",
x"7AC46817",
x"7AEA6831",
x"7B176834",
x"7B53681B",
x"7BA567EB",
x"7C0E67A7",
x"7C936758",
x"7D326707",
x"7DEA66C2",
x"7EB56690",
x"7F8C6679",
x"80626681",
x"812A66AA",
x"81D866EC",
x"825D673E",
x"82B16799",
x"82CB67ED",
x"82A76832",
x"82486860",
x"81B76873",
x"80FD6868",
x"802B6842",
x"7F4F6807",
x"7E7A67BE",
x"7DBA676D",
x"7D19671D",
x"7C9B66D2",
x"7C46668E",
x"7C196658",
x"7C0D662E",
x"7C1A660D",
x"7C3865F7",
x"7C5C65E8",
x"7C7F65DB",
x"7C9465D0",
x"7C9765C5",
x"7C8465B7",
x"7C5965A4",
x"7C14658D",
x"7BBC6572",
x"7B536555",
x"7AE36538",
x"7A72651D",
x"7A096509",
x"79AE64FD",
x"796964FA",
x"793F6504",
x"79306517",
x"793B6535",
x"795F655B",
x"79966586",
x"79D865B5",
x"7A2065E3",
x"7A69660E",
x"7AAE6635",
x"7AEF6655",
x"7B2B666A",
x"7B666675",
x"7BA36673",
x"7BE36660",
x"7C28663C",
x"7C6F6601",
x"7CAA65AF",
x"7CCC653F",
x"7CBE64AE",
x"7C6563F7",
x"7BA16318",
x"7A59620A",
x"787760CC",
x"75F05F5D",
x"72C85DC2",
x"6F135BFE",
x"6AF95A1F",
x"66B15838",
x"627D565C",
x"5EA754A6",
x"5B785335",
x"592D5222",
x"57F65189",
x"57EF517C",
x"59195204",
x"5B5B531C",
x"5E8A54BA",
x"626956C3",
x"66B15917",
x"6B195B8D",
x"6F5E5E01",
x"7348604F",
x"76AE625A",
x"79796413",
x"7BA1656F",
x"7D2E6672",
x"7E326725",
x"7EC5679A",
x"7F0167E2",
x"7F01680A",
x"7ED96820",
x"7E9E682A",
x"7E5F682D",
x"7E256826",
x"7DF96814",
x"7DE067F9",
x"7DDF67D3",
x"7DF767AB",
x"7E276783",
x"7E6C6766",
x"7EC1675C",
x"7F20676B",
x"7F806793",
x"7FD967D2",
x"80256826",
x"805D6880",
x"807E68D9",
x"808A6926",
x"8083695F",
x"806C6982",
x"804B698E",
x"8027698A",
x"8006697F",
x"7FEA6975",
x"7FD96977",
x"7FD3698C",
x"7FDB69BA",
x"7FF069FF",
x"80186A5B",
x"80536AC9",
x"80A56B42",
x"810E6BBE",
x"81916C37",
x"822D6CA4",
x"82DC6D03",
x"83986D4E",
x"84566D80",
x"850A6D97",
x"85A86D92",
x"86256D6B",
x"86766D27",
x"869A6CC7",
x"86916C52",
x"86656BD2",
x"86216B52",
x"85D96AE2",
x"85A06A8F",
x"85876A63",
x"85A16A6B",
x"85F66AA7",
x"86866B13",
x"87486BA7",
x"882E6C52",
x"89226D02",
x"8A096DA1",
x"8AC66E20",
x"8B446E6F",
x"8B716E89",
x"8B456E6F",
x"8ABF6E27",
x"89EA6DBE",
x"88D86D44",
x"879E6CC5",
x"86556C4F",
x"85116BE6",
x"83E56B89",
x"82DA6B32",
x"81F66AD9",
x"81356A70",
x"809369EF",
x"8007694F",
x"7F8D6894",
x"7F1B67C2",
x"7EB566E9",
x"7E596617",
x"7E0B6560",
x"7DD364CF",
x"7DB26470",
x"7DAB6444",
x"7DB86445",
x"7DD36468",
x"7DF5649D",
x"7E0D64D6",
x"7E136504",
x"7DFF6520",
x"7DCC6525",
x"7D84651B",
x"7D31650D",
x"7CE36507",
x"7CAF651B",
x"7CAD6552",
x"7CEA65B7",
x"7D726648",
x"7E416700",
x"7F4B67D2",
x"807968A8",
x"81A5696F",
x"82AB6A0D",
x"83606A6F",
x"83A16A86",
x"83566A47",
x"827669B2",
x"810668D4",
x"7F2267BC",
x"7CF46684",
x"7AB4654E",
x"78A06438",
x"76F9636A",
x"75F76301",
x"75CF6317",
x"769D63BC",
x"786F64F7",
x"7B3F66C2",
x"7EF6690C",
x"836A6BB8",
x"886A6EA7",
x"8DB871B3",
x"931A74B7",
x"98597796",
x"9D487A34",
x"A1C27C86",
x"A5B97E87",
x"A928803A",
x"AC1981B2",
x"AEA682FE",
x"B0EE8433",
x"B3148566",
x"B535869F",
x"B76A87E7",
x"B9C0893B",
x"BC388A91",
x"BEC38BDA",
x"C14D8D03",
x"C3B78DF9",
x"C5E48EAC",
x"C7B98F14",
x"C9238F2C",
x"CA1D8EFD",
x"CAB28E91",
x"CAF18DFD",
x"CAFB8D56",
x"CAEF8CB8",
x"CAEF8C35",
x"CB198BE3",
x"CB7E8BCF",
x"CC288C03",
x"CD128C7D",
x"CE338D3E",
x"CF7B8E3C",
x"D0D88F6D",
x"D23990C5",
x"D3959235",
x"D4E493AF",
x"D6299527",
x"D76B9691",
x"D8B397E5",
x"DA0B991A",
x"DB799A2D",
x"DD029B1A",
x"DEA29BE2",
x"E0509C86",
x"E1FB9D09",
x"E3929D71",
x"E4FC9DBD",
x"E6249DEF",
x"E6F69E08",
x"E7629E05",
x"E75F9DDE",
x"E6EB9D93",
x"E6099D1D",
x"E4CA9C7D",
x"E3419BB8",
x"E1899AD7",
x"DFC499E5",
x"DE0D98FB",
x"DC88982B",
x"DB48978C",
x"DA61972D",
x"D9DA971D",
x"D9B3975B",
x"D9DF97E4",
x"DA5098A4",
x"DAE8998A",
x"DB939A7B",
x"DC339B5A",
x"DCB19C0F",
x"DCFE9C89",
x"DD0B9CBD",
x"DCD19CA7",
x"DC579C52",
x"DBA59BCC",
x"DAC99B27",
x"D9D59A79",
x"D8E299D8",
x"D809995A",
x"D75D990A",
x"D6F198F2",
x"D6D19914",
x"D703996C",
x"D78299EE",
x"D8439A8A",
x"D92E9B31",
x"DA2F9BD2",
x"DB299C5B",
x"DC039CC1",
x"DCAC9CFD",
x"DD179D10",
x"DD489D00",
x"DD449CDB",
x"DD1D9CB0",
x"DCE79C8D",
x"DCB49C82",
x"DC969C9A",
x"DC929CD5",
x"DCA69D33",
x"DCCA9DA4",
x"DCEB9E1C",
x"DCF99E83",
x"DCE59ECD",
x"DCA69EE8",
x"DC3B9ED0",
x"DBB39E82",
x"DB199E08",
x"DA809D6C",
x"D9F99CBB",
x"D9859BFF",
x"D9159B3B",
x"D88C9A69",
x"D7B79979",
x"D65B9856",
x"D43696E2",
x"D10C9503",
x"CCB292A0",
x"C7188FAE",
x"C04D8C31",
x"B884883B",
x"B00E83EE",
x"A7547F7B",
x"9ECC7B18",
x"96EA76FC",
x"9018735F",
x"8AA8706B",
x"86CF6E3B",
x"84A16CDE",
x"84156C54",
x"85096C8A",
x"874B6D6C",
x"8A9E6ED9",
x"8EC870B1",
x"938E72D7",
x"98BF752F",
x"9E3277A0",
x"A3C27A1B",
x"A9507C8F",
x"AEBC7EF1",
x"B3EB8136",
x"B8BF835A",
x"BD1C8554",
x"C0ED8721",
x"C42288BB",
x"C6B78A22",
x"C8B38B5A",
x"CA288C67",
x"CB2D8D4C",
x"CBE18E10",
x"CC608EB8",
x"CCC18F4B",
x"CD198FC8",
x"CD6F9037",
x"CDC69094",
x"CE1890E5",
x"CE60912A",
x"CE969169",
x"CEB991A5",
x"CEC991E3",
x"CECB922A",
x"CEC7927A",
x"CEC392D6",
x"CEC3933A",
x"CEC1939E",
x"CEB993F9",
x"CE9C943F",
x"CE589465",
x"CDE09462",
x"CD27942E",
x"CC2C93CC",
x"CAF89344",
x"C9A0929D",
x"C84691EC",
x"C70E9142",
x"C62590B5",
x"C5B09055",
x"C5D1902F",
x"C6999049",
x"C80890A4",
x"CA0F9135",
x"CC8B91F3",
x"CF4E92C9",
x"D22393A8",
x"D4CE947D",
x"D71C953A",
x"D8E195D2",
x"DA009641",
x"DA6E968A",
x"DA3496B0",
x"D96996BD",
x"D83796BD",
x"D6C896B8",
x"D55396BA",
x"D40296C7",
x"D2FE96E4",
x"D25D9710",
x"D22A974A",
x"D267978C",
x"D30197D2",
x"D3E4981B",
x"D4F59865",
x"D61C98B0",
x"D74398FB",
x"D85A9948",
x"D958999A",
x"DA3B99EE",
x"DB029A3D",
x"DBB09A83",
x"DC479AB4",
x"DCC39AC5",
x"DD219AAD",
x"DD5B9A64",
x"DD6B99E4",
x"DD4A9933",
x"DCF5985B",
x"DC6F976E",
x"DBC09682",
x"DAF595AE",
x"DA1C950D",
x"D94794AF",
x"D88394A0",
x"D7DA94E0",
x"D74A9568",
x"D6D0961E",
x"D66096EB",
x"D5E497AA",
x"D54B983A",
x"D47E987C",
x"D36B9859",
x"D20697C7",
x"D04A96C2",
x"CE399555",
x"CBDD9394",
x"C942919B",
x"C67F8F87",
x"C3A88D7A",
x"C0D48B90",
x"BE1989DF",
x"BB878877",
x"B928875D",
x"B6FD868F",
x"B4FE85FD",
x"B3188591",
x"B12D852E",
x"AF1484AC",
x"AC9B83E8",
x"A98E82B9",
x"A5BF8100",
x"A1057EA2",
x"9B507B93",
x"94A277DA",
x"8D1D738B",
x"84FF6ECE",
x"7C9B69D8",
x"745F64EC",
x"6CBB604D",
x"661E5C3F",
x"60E858F5",
x"5D5C569C",
x"5B9C5543",
x"5BA154E7",
x"5D415570",
x"603156B6",
x"64135884",
x"687C5AA4",
x"6D075CDF",
x"715C5F0B",
x"75376107",
x"786F62C4",
x"7AF96439",
x"7CDE656F",
x"7E3A6672",
x"7F356752",
x"7FFD681D",
x"80B868E1",
x"818769A6",
x"827E6A6D",
x"83AB6B3B",
x"850A6C0D",
x"86946CE1",
x"88386DB7",
x"89E26E8F",
x"8B806F68",
x"8D007043",
x"8E52711F",
x"8F6E71F6",
x"905072C4",
x"90F9737F",
x"91707420",
x"91C2749C",
x"91FD74EC",
x"9231750D",
x"926C7502",
x"92B974D1",
x"93227483",
x"93A8742A",
x"944973DA",
x"950173A5",
x"95C9739C",
x"969A73D0",
x"9770744A",
x"984A750D",
x"992E7615",
x"9A1C7754",
x"9B2178BA",
x"9C427A30",
x"9D847B9C",
x"9EE77CE5",
x"A0637DFA",
x"A1ED7EC7",
x"A3717F49",
x"A4DC7F81",
x"A6177F7A",
x"A7117F42",
x"A7C07EF1",
x"A8257E9C",
x"A84A7E5A",
x"A8477E40",
x"A83F7E5D",
x"A8577EBA",
x"A8BF7F60",
x"A99C8050",
x"AB11818A",
x"AD308304",
x"B00184BC",
x"B37286A2",
x"B76388AC",
x"BBA38AC8",
x"BFF88CDF",
x"C41C8EDF",
x"C7D090AF",
x"CAD7923D",
x"CD059376",
x"CE40944E",
x"CE8194C5",
x"CDD894DE",
x"CC6A94A4",
x"CA6B942D",
x"C819938D",
x"C5B392D8",
x"C3759221",
x"C1919174",
x"C02590DC",
x"BF3D9055",
x"BED48FDC",
x"BED18F69",
x"BF0F8EF3",
x"BF608E71",
x"BF988DDF",
x"BF918D39",
x"BF308C83",
x"BE6D8BBE",
x"BD508AF4",
x"BBEE8A2C",
x"BA6A8971",
x"B8F188C9",
x"B7AB8840",
x"B6C087DD",
x"B64A87A7",
x"B65487A1",
x"B6DA87D0",
x"B7C7882F",
x"B8FB88BB",
x"BA498964",
x"BB878A1D",
x"BC8B8ACF",
x"BD328B67",
x"BD658BD2",
x"BD1C8BFB",
x"BC548BDA",
x"BB198B69",
x"B9748AA5",
x"B7748995",
x"B51F883F",
x"B27886A8",
x"AF7884D6",
x"AC1582CA",
x"A83F8082",
x"A3F07DFE",
x"9F287B3A",
x"99F7783C",
x"947E7510",
x"8EF071CE",
x"898D6E93",
x"849B6B87",
x"806368D5",
x"7D2166A3",
x"7B036513",
x"7A186438",
x"7A5B6415",
x"7BAA64A0",
x"7DCF65BC",
x"80876744",
x"83906910",
x"86AB6AF6",
x"89A96CD9",
x"8C716EA3",
x"8EFD704D",
x"915671DF",
x"9398736A",
x"95E274FF",
x"985076B6",
x"9AFB789B",
x"9DEC7AB6",
x"A11F7D01",
x"A4887F6D",
x"A80D81E7",
x"AB918453",
x"AEF78699",
x"B22C88A4",
x"B5198A62",
x"B7B78BCC",
x"BA028CE0",
x"BBF88DA4",
x"BD9F8E20",
x"BEFA8E60",
x"C00F8E6F",
x"C0E08E56",
x"C1718E1D",
x"C1CA8DCE",
x"C1F28D6F",
x"C1F48D0B",
x"C1E38CB1",
x"C1D08C6D",
x"C1D38C53",
x"C2018C74",
x"C26F8CE0",
x"C32A8DA2",
x"C43C8EC1",
x"C5A39038",
x"C75A91FC",
x"C95093F6",
x"CB729609",
x"CDA99817",
x"CFDD99FD",
x"D1F79B9F",
x"D3E79CE8",
x"D5A29DCD",
x"D7239E4B",
x"D8699E73",
x"D97B9E55",
x"DA5A9E0F",
x"DB0B9DB7",
x"DB939D69",
x"DBF19D33",
x"DC209D19",
x"DC1D9D16",
x"DBE79D1C",
x"DB7E9D15",
x"DAEA9CE5",
x"DA3A9C79",
x"D9869BC1",
x"D8E59AB7",
x"D873995F",
x"D84697CA",
x"D867960A",
x"D8D5943E",
x"D982927D",
x"DA5190DC",
x"DB198F69",
x"DBB08E2B",
x"DBEF8D24",
x"DBBB8C4F",
x"DB068BA8",
x"D9D78B2A",
x"D8468AD3",
x"D6788AA8",
x"D49C8AAC",
x"D2DF8AE7",
x"D1658B5A",
x"D0408C04",
x"CF728CDA",
x"CEE78DC9",
x"CE788EB7",
x"CDF28F81",
x"CD259009",
x"CBDD902D",
x"C9F88FD6",
x"C7648EFA",
x"C4258D97",
x"C0538BBE",
x"BC188985",
x"B7AB8714",
x"B34A8492",
x"AF338229",
x"AB9E7FFE",
x"A8AC7E33",
x"A6787CD9",
x"A5047BF7",
x"A43F7B89",
x"A4047B7F",
x"A4227BBD",
x"A4607C22",
x"A4827C85",
x"A4527CC4",
x"A3A57CC0",
x"A2637C61",
x"A0857B9E",
x"9E1C7A75",
x"9B4C78F7",
x"9840773C",
x"952F7564",
x"924C7390",
x"8FBE71E2",
x"8D9B706F",
x"8BE66F45",
x"8A8D6E65",
x"896A6DBE",
x"88526D3D",
x"87116CC1",
x"857B6C2D",
x"83766B66",
x"80F66A5F",
x"7E0B6911",
x"7ADC6786",
x"779A65D3",
x"74866418",
x"71DC627A",
x"6FD6611A",
x"6E9B6015",
x"6E3F5F84",
x"6EC25F70",
x"70105FD6",
x"720660AD",
x"747461DC",
x"7731634F",
x"7A0D64EC",
x"7CE9669A",
x"7FAA6848",
x"824369E5",
x"84B56B6B",
x"86FD6CD4",
x"89246E21",
x"8B2E6F57",
x"8D1D7076",
x"8EF07183",
x"90A17285",
x"9228737C",
x"937E746C",
x"949C7557",
x"9581763A",
x"96337718",
x"96BC77E8",
x"972B78A7",
x"9791794E",
x"980179D4",
x"988A7A33",
x"99367A67",
x"9A0A7A72",
x"9B057A5D",
x"9C1F7A33",
x"9D507A09",
x"9E8879F4",
x"9FBF7A08",
x"A0EB7A58",
x"A2087AF1",
x"A3177BD3",
x"A41C7CFB",
x"A5217E5B",
x"A62F7FDB",
x"A74F8168",
x"A88B82E7",
x"A9E68445",
x"AB5E8571",
x"ACF38666",
x"AE95871F",
x"B03F87A2",
x"B1DD87F4",
x"B363881D",
x"B4BF8822",
x"B5E38808",
x"B6C287D3",
x"B7518783",
x"B78E8717",
x"B774868E",
x"B70A85EC",
x"B6578533",
x"B56E846C",
x"B45E839F",
x"B34482D7",
x"B236821F",
x"B1518185",
x"B0AF8111",
x"B06480CF",
x"B08180C7",
x"B10B80FE",
x"B2048178",
x"B35D8230",
x"B5058321",
x"B6DE843C",
x"B8CA8571",
x"BAA386A8",
x"BC4987C8",
x"BDA088B9",
x"BE948969",
x"BF1889CA",
x"BF2D89DC",
x"BEE089A1",
x"BE43892B",
x"BD71888E",
x"BC8887E6",
x"BBA38748",
x"BADE86C9",
x"BA4A8677",
x"B9F28653",
x"B9D98659",
x"B9F7867E",
x"BA4086B3",
x"BAA586E6",
x"BB0F8707",
x"BB70870E",
x"BBB386F3",
x"BBCD86B6",
x"BBB6865D",
x"BB6A85EC",
x"BAED856C",
x"BA4684E6",
x"B9828466",
x"B8AF83F1",
x"B7DE8392",
x"B720834F",
x"B682832D",
x"B60E8333",
x"B5C4835C",
x"B5A683A6",
x"B5A68408",
x"B5B68474",
x"B5C984DE",
x"B5CD8538",
x"B5BC8577",
x"B5918598",
x"B5508599",
x"B5048587",
x"B4BA8568",
x"B47B854C",
x"B4468535",
x"B4118523",
x"B3BD850B",
x"B32184D3",
x"B2018457",
x"B0248372",
x"AD508200",
x"A9607FE3",
x"A4427D11",
x"9E077990",
x"96E67582",
x"8F31711A",
x"87586C9A",
x"7FD2684E",
x"791A647C",
x"73976160",
x"6F995F25",
x"6D445DDA",
x"6C9B5D7A",
x"6D785DE9",
x"6F945EF8",
x"72966072",
x"7619621D",
x"79C163C8",
x"7D3C654C",
x"804F6690",
x"82D8678C",
x"84C96842",
x"862F68C2",
x"871E691D",
x"87B76968",
x"881869B2",
x"88606A09",
x"88A46A6F",
x"88EF6AE5",
x"89466B61",
x"89A96BD9",
x"8A106C44",
x"8A736C9A",
x"8AC96CD7",
x"8B116CF9",
x"8B456D08",
x"8B696D0C",
x"8B7F6D0C",
x"8B8B6D14",
x"8B946D2A",
x"8B9D6D54",
x"8BA76D8D",
x"8BAF6DD2",
x"8BB26E1A",
x"8BAA6E5C",
x"8B8E6E8C",
x"8B586EA1",
x"8B016E96",
x"8A8B6E68",
x"89FC6E1A",
x"89596DB1",
x"88B46D38",
x"881D6CB7",
x"87A76C3A",
x"87626BCC",
x"875D6B78",
x"87A06B44",
x"88286B35",
x"88F06B4F",
x"89E96B93",
x"8B046BFD",
x"8C2B6C89",
x"8D4F6D2D",
x"8E606DDF",
x"8F586E94",
x"902F6F43",
x"90ED6FDB",
x"91947057",
x"922970AD",
x"92B570D8",
x"933470DA",
x"93A270AD",
x"93F6705A",
x"94206FDF",
x"94106F45",
x"93B86E92",
x"93106DC8",
x"92156CF3",
x"90D66C1C",
x"8F666B4E",
x"8DE36A97",
x"8C736A06",
x"8B3B69A8",
x"8A5D698C",
x"89F069B5",
x"8A036A27",
x"8A916ADC",
x"8B8A6BC5",
x"8CCF6CCF",
x"8E3C6DE6",
x"8FA86EF0",
x"90ED6FD9",
x"91EC7093",
x"92907116",
x"92D2715F",
x"92B57178",
x"9249716B",
x"91A27147",
x"90D8711A",
x"900170F2",
x"8F3270D5",
x"8E7970C7",
x"8DDB70C7",
x"8D5C70CF",
x"8CFA70DB",
x"8CB470E4",
x"8C8170E5",
x"8C6370DE",
x"8C5670D1",
x"8C5C70BE",
x"8C7770AB",
x"8CA5709C",
x"8CE77093",
x"8D3B708D",
x"8D97708D",
x"8DF6708D",
x"8E4C708A",
x"8E927080",
x"8EBC706B",
x"8EC57048",
x"8EA47017",
x"8E576FD7",
x"8DDC6F83",
x"8D2E6F1A",
x"8C4B6E96",
x"8B2B6DF0",
x"89C96D21",
x"88206C20",
x"86276AE8",
x"83DA6975",
x"814167CC",
x"7E5F65F7",
x"7B496407",
x"78186213",
x"74EF6033",
x"71F05E87",
x"6F425D25",
x"6D075C21",
x"6B5C5B88",
x"6A4E5B5C",
x"69E15B97",
x"6A0F5C25",
x"6AC45CF1",
x"6BE55DE3",
x"6D545EDD",
x"6EF05FCC",
x"70A3609F",
x"72526150",
x"73F661E0",
x"7589625A",
x"770D62CC",
x"788C6345",
x"7A0E63D6",
x"7BA1648D",
x"7D4B656D",
x"7F0E6679",
x"80ED67A7",
x"82E368EF",
x"84E66A42",
x"86EA6B90",
x"88E26CCD",
x"8ABE6DEC",
x"8C736EE6",
x"8DF46FBA",
x"8F397066",
x"904170EE",
x"91067154",
x"918E719D",
x"91E371CF",
x"920B71EE",
x"921471FE",
x"92097202",
x"91F47200",
x"91E071FB",
x"91D371F6",
x"91CF71F4",
x"91D571F4",
x"91E071F8",
x"91F071FE",
x"92037203",
x"92157209",
x"922E7210",
x"924E721C",
x"92807231",
x"92C97258",
x"93357299",
x"93C572FB",
x"947E7383",
x"955D7430",
x"965D74FC",
x"977675DB",
x"989A76BC",
x"99BF778B",
x"9ADA7833",
x"9BE378A7",
x"9CD278DE",
x"9DA178D6",
x"9E507893",
x"9EDD7829",
x"9F4977AC",
x"9F947733",
x"9FBF76D5",
x"9FCD76A6",
x"9FC576AF",
x"9FAC76F4",
x"9F8B7771",
x"9F6E7816",
x"9F6078D4",
x"9F6C7993",
x"9F987A40",
x"9FE97AC9",
x"A05D7B22",
x"A0ED7B43",
x"A18A7B2D",
x"A2257AE7",
x"A2A97A7B",
x"A30879F4",
x"A32F7961",
x"A31778CE",
x"A2BB7844",
x"A21C77CB",
x"A1457765",
x"A03E7710",
x"9F1476CA",
x"9DD7768B",
x"9C91764A",
x"9B4B7601",
x"9A0575A5",
x"98C5752F",
x"9784749A",
x"964273E2",
x"94F97309",
x"93A87210",
x"924E70FC",
x"90EE6FD8",
x"8F8E6EAD",
x"8E366D89",
x"8CF06C7C",
x"8BC26B96",
x"8AB66ADF",
x"89D26A66",
x"89146A2B",
x"887C6A31",
x"88046A6D",
x"87A46AD5",
x"87536B59",
x"87076BE5",
x"86B86C66",
x"865F6CCE",
x"85F96D0F",
x"85816D1E",
x"84F66CFC",
x"84536CAB",
x"83956C2E",
x"82B96B8D",
x"81B56ACF",
x"808369F9",
x"7F1D6911",
x"7D806819",
x"7BB26711",
x"79BF6601",
x"77BA64EC",
x"75BA63D8",
x"73DF62CF",
x"724861DC",
x"7111610D",
x"704C606A",
x"70055FFE",
x"70355FC9",
x"70D45FCD",
x"71C86006",
x"72F76069",
x"744760F0",
x"759D6190",
x"76EF6243",
x"78376309",
x"797C63DF",
x"7AD164CB",
x"7C4665D0",
x"7DF366F6",
x"7FE7683B",
x"822B69A1",
x"84BE6B21",
x"87906CB1",
x"8A8E6E45",
x"8D9C6FD1",
x"909D7147",
x"9374729D",
x"960B73CE",
x"985674D7",
x"9A4D75BD",
x"9BF17683",
x"9D4C7734",
x"9E6677D5",
x"9F4D786D",
x"A00B78FB",
x"A0A97981",
x"A12F79F9",
x"A19C7A5E",
x"A1F17AAA",
x"A2307AD7",
x"A2567ADE",
x"A2667ABE",
x"A2617A7B",
x"A24F7A18",
x"A2357999",
x"A221790C",
x"A21E7879",
x"A23C77EE",
x"A28A7777",
x"A3147720",
x"A3E676F4",
x"A50476FB",
x"A66D773A",
x"A81777B4",
x"A9ED7867",
x"ABD77948",
x"ADB57A4D",
x"AF647B64",
x"B0C57C7E",
x"B1B97D85",
x"B2327E68",
x"B2287F1B",
x"B1A17F96",
x"B0B07FD9",
x"AF737FE4",
x"AE0D7FC3",
x"ACA27F82",
x"AB527F2D",
x"AA3B7ED3",
x"A96D7E7A",
x"A8F37E29",
x"A8CD7DE5",
x"A8F37DB0",
x"A9567D85",
x"A9EA7D65",
x"AA9E7D4E",
x"AB5E7D41",
x"AC1F7D3F",
x"ACD27D47",
x"AD647D5D",
x"ADD27D7C",
x"AE0B7DA5",
x"AE0B7DCF",
x"ADCD7DF1",
x"AD547E04",
x"ACAD7E01",
x"ABE47DE5",
x"AB127DB3",
x"AA517D72",
x"A9BF7D30",
x"A9707CFE",
x"A9737CE8",
x"A9C97CFB",
x"AA667D3C",
x"AB317DA3",
x"AC047E28",
x"ACB37EAD",
x"AD117F19",
x"ACF47F53",
x"AC427F3C",
x"AAEB7EC9",
x"A8F57DED",
x"A6777CB2",
x"A3927B29",
x"A07A796E",
x"9D6077A3",
x"9A7775E7",
x"97E77458",
x"95CC730B",
x"9434720A",
x"931A7158",
x"926C70E9",
x"920D70B1",
x"91DA709A",
x"91AF7092",
x"91707085",
x"91017068",
x"90597034",
x"8F776FE4",
x"8E636F79",
x"8D2C6EF9",
x"8BE66E65",
x"8A9F6DC2",
x"89666D10",
x"88386C4E",
x"87106B76",
x"85DB6A84",
x"84816975",
x"82EC6844",
x"810166F2",
x"7EB56584",
x"7C096407",
x"79096286",
x"75D56115",
x"72975FC8",
x"6F855EAF",
x"6CD15DDA",
x"6AB05D55",
x"69455D1E",
x"68A45D33",
x"68D25D88",
x"69BA5E0A",
x"6B385EA7",
x"6D1E5F46",
x"6F375FD6",
x"714E604B",
x"73376098",
x"74CF60C1",
x"760760C8",
x"76DC60BB",
x"775B60A8",
x"779B60A1",
x"77BF60B5",
x"77E660F3",
x"78326163",
x"78BA6209",
x"798E62E2",
x"7AB763E5",
x"7C2D6506",
x"7DE06637",
x"7FBF6763",
x"81AB687D",
x"838D6973",
x"85486A3D",
x"86C96AD2",
x"88036B37",
x"88F26B6D",
x"899A6B86",
x"8A076B8D",
x"8A4C6B96",
x"8A816BAD",
x"8ABB6BDE",
x"8B116C31",
x"8B936CA6",
x"8C496D37",
x"8D386DDB",
x"8E596E85",
x"8FA56F29",
x"910B6FBE",
x"927E7043",
x"93ED70B5",
x"954D7121",
x"96977192",
x"97C87216",
x"98E372BA",
x"99EF7389",
x"9AF67485",
x"9C0075AA",
x"9D1576EE",
x"9E3B7840",
x"9F6D7989",
x"A0A57AB7",
x"A1D57BB4",
x"A2EE7C75",
x"A3DC7CEF",
x"A48D7D26",
x"A4F47D1C",
x"A5077CE0",
x"A4C77C7F",
x"A43C7C0C",
x"A3737B93",
x"A2847B23",
x"A1857AC6",
x"A0917A7C",
x"9FBB7A4B",
x"9F127A2C",
x"9E9E7A19",
x"9E607A0C",
x"9E4F79F9",
x"9E6079DA",
x"9E8779AA",
x"9EB67965",
x"9EE6790C",
x"9F1178A5",
x"9F3B7834",
x"9F6777C7",
x"9F9E7765",
x"9FE77718",
x"A04876E7",
x"A0C276D2",
x"A15076DA",
x"A1EA76F4",
x"A2857716",
x"A3117733",
x"A37D773A",
x"A3BB7723",
x"A3BF76E1",
x"A3807675",
x"A2F775E2",
x"A224752F",
x"A1077468",
x"9FA7739C",
x"9E0A72D8",
x"9C3C7227",
x"9A4D7190",
x"98507116",
x"965770B9",
x"94797073",
x"92C67041",
x"9153701C",
x"90286FFE",
x"8F466FDF",
x"8EA86FC1",
x"8E416F9C",
x"8DFD6F6C",
x"8DC86F30",
x"8D8D6EE4",
x"8D3E6E83",
x"8CD66E0C",
x"8C556D80",
x"8BC66CE2",
x"8B356C37",
x"8AB16B87",
x"8A426ADE",
x"89E96A41",
x"899B69B8",
x"89436944",
x"88BF68E1",
x"87EC6883",
x"86A7681B",
x"84D26799",
x"826366E6",
x"7F5B65F9",
x"7BD264C8",
x"77F26356",
x"73F061AE",
x"70095FE3",
x"6C7C5E10",
x"697D5C52",
x"67375AC7",
x"65C15988",
x"652458A9",
x"65555832",
x"663D5824",
x"67BD5878",
x"69B05924",
x"6BF65A17",
x"6E6D5B3F",
x"70FD5C90",
x"73965DFE",
x"76275F84",
x"78AD611A",
x"7B2162BE",
x"7D83646A",
x"7FD2661E",
x"821067CF",
x"84396975",
x"86526B06",
x"88596C75",
x"8A506DBB",
x"8C396ED2",
x"8E156FB9",
x"8FE37072",
x"91A47109",
x"9355718A",
x"94F37205",
x"967A7286",
x"97E6731A",
x"993273C8",
x"9A5C7492",
x"9B617572",
x"9C407660",
x"9CF8774B",
x"9D8D7827",
x"9DFD78E2",
x"9E4D7972",
x"9E8379CB",
x"9E9F79ED",
x"9EAC79D7",
x"9EB27995",
x"9EBB7933",
x"9ED378C1",
x"9F0B7854",
x"9F7477FB",
x"A01B77C8",
x"A10D77C6",
x"A24D77FB",
x"A3DF7865",
x"A5B678FF",
x"A7C279BE",
x"A9E97A93",
x"AC0B7B6B",
x"AE077C36",
x"AFC07CE5",
x"B11E7D6F",
x"B20E7DCF",
x"B28C7E02",
x"B2A37E0F",
x"B2647DFE",
x"B1EB7DD9",
x"B15A7DAA",
x"B0D37D7F",
x"B0717D60",
x"B0507D51",
x"B07A7D5B",
x"B0F47D7E",
x"B1B97DC0",
x"B2BF7E1F",
x"B3F37EA0",
x"B5447F43",
x"B6A5800C",
x"B80880F8",
x"B9678207",
x"BABC832D",
x"BBFF8464",
x"BD32859C",
x"BE4986C5",
x"BF3A87CA",
x"BFFC889D",
x"C07F8929",
x"C0B38969",
x"C08F8958",
x"C00988F7",
x"BF238853",
x"BDE4877E",
x"BC5B868A",
x"BA9B858E",
x"B8B9849F",
x"B6CD83D0",
x"B4ED832B",
x"B32682B8",
x"B1878272",
x"B0148257",
x"AED08257",
x"ADBA8266",
x"ACD38271",
x"AC14826A",
x"AB7E8246",
x"AB0C81FB",
x"AAB98185",
x"AA7E80E4",
x"AA50801B",
x"AA1E7F2F",
x"A9D67E2A",
x"A9677D11",
x"A8BF7BEF",
x"A7D37AD3",
x"A6A179C3",
x"A52B78CA",
x"A38177F2",
x"A1B87741",
x"9FEA76BC",
x"9E2E765E",
x"9C987623",
x"9B3175FB",
x"99F775D5",
x"98DA759A",
x"97C27537",
x"968D7495",
x"951A73A7",
x"9350726A",
x"911F70DF",
x"8E876F1C",
x"8B9B6D3A",
x"887E6B59",
x"855C69A3",
x"826D6837",
x"7FE26731",
x"7DE966A1",
x"7C9E668B",
x"7C1366E5",
x"7C416796",
x"7D196883",
x"7E7F698A",
x"80536A90",
x"827A6B7F",
x"84DA6C4E",
x"87666D00",
x"8A156DA3",
x"8CEC6E4D",
x"8FED6F19",
x"9321701F",
x"96867170",
x"9A177319",
x"9DC67512",
x"A17E774B",
x"A52279AD",
x"A8957C15",
x"ABBC7E63",
x"AE7E8074",
x"B0CD8233",
x"B2A68392",
x"B40C848D",
x"B50E8529",
x"B5BF8578",
x"B6388592",
x"B68F858E",
x"B6DB8585",
x"B72D858A",
x"B78F85A9",
x"B80485EA",
x"B88A864A",
x"B91986C5",
x"B9A9874F",
x"BA2F87DF",
x"BAA3886A",
x"BAFF88EA",
x"BB478960",
x"BB7E89D0",
x"BBB08A3F",
x"BBEB8AB9",
x"BC3C8B46",
x"BCB28BEF",
x"BD598CB6",
x"BE358D9D",
x"BF498E9E",
x"C0928FB1",
x"C20790CB",
x"C39E91DF",
x"C54692E2",
x"C6F493CB",
x"C8959494",
x"CA19953A",
x"CB6F95BB",
x"CC829616",
x"CD3F964C",
x"CD95965B",
x"CD729641",
x"CCD195FC",
x"CBB0958A",
x"CA1D94EC",
x"C8339425",
x"C6169341",
x"C3F7924B",
x"C2089155",
x"C07F9073",
x"BF848FB9",
x"BF328F3C",
x"BF928F07",
x"C0988F22",
x"C2268F8E",
x"C40E9042",
x"C6189132",
x"C80E924C",
x"C9BD9379",
x"CB0294A1",
x"CBC795B1",
x"CC069693",
x"CBCA9735",
x"CB23978D",
x"CA2C978C",
x"C8F99730",
x"C7A09675",
x"C628955C",
x"C49493F0",
x"C2DE923D",
x"C101904E",
x"BEF28E3B",
x"BCAF8C17",
x"BA3989F9",
x"B79887F3",
x"B4DC8617",
x"B219846E",
x"AF6B8300",
x"ACE881CA",
x"AAA380C9",
x"A8AC7FF4",
x"A70B7F40",
x"A5C27EA6",
x"A4CA7E1C",
x"A41A7D9E",
x"A3A27D26",
x"A3527CB6",
x"A3187C50",
x"A2E77BF5",
x"A2B37BA8",
x"A2767B67",
x"A22E7B36",
x"A1DF7B15",
x"A1947AFF",
x"A1597AF8",
x"A13B7AFC",
x"A1427B0B",
x"A1717B1C",
x"A1BE7B2C",
x"A20E7B2A",
x"A23C7B06",
x"A2107AAA",
x"A14A79FC",
x"9FAF78E4",
x"9D06774D",
x"992C752A",
x"9418727E",
x"8DE76F57",
x"86D56BD7",
x"7F44682A",
x"77A8648A",
x"708C6134",
x"6A6C5E5F",
x"65BD5C3B",
x"62CA5AE7",
x"61C05A70",
x"62975ACC",
x"65285BE3",
x"69235D8E",
x"6E245F9F",
x"73C861EA",
x"79A86448",
x"7F776699",
x"84FB68CE",
x"8A156ADE",
x"8EBC6CCF",
x"92F66EA9",
x"96D27073",
x"9A5F7234",
x"9DA473EB",
x"A09E7592",
x"A33D771D",
x"A573787C",
x"A72479A0",
x"A8407A81",
x"A8C27B19",
x"A8AE7B6D",
x"A8197B86",
x"A72B7B78",
x"A60A7B57",
x"A4E37B37",
x"A3E17B28",
x"A3247B33",
x"A2B87B5A",
x"A29E7B99",
x"A2C77BE1",
x"A3187C28",
x"A36D7C5A",
x"A3A27C6D",
x"A39F7C59",
x"A34D7C1E",
x"A2AC7BC3",
x"A1C67B54",
x"A0AF7AE4",
x"9F8B7A82",
x"9E7E7A41",
x"9DAB7A2D",
x"9D2C7A49",
x"9D157A92",
x"9D6A7AFE",
x"9E1F7B7E",
x"9F1F7BFC",
x"A04D7C65",
x"A1857CA6",
x"A2A87CAF",
x"A39B7C7E",
x"A44F7C11",
x"A4BC7B74",
x"A4E77AB9",
x"A4DE79F2",
x"A4B17939",
x"A471789F",
x"A42C7833",
x"A3E977FB",
x"A3A577F4",
x"A3567812",
x"A2EE7846",
x"A25F7879",
x"A19A7899",
x"A09B7895",
x"9F697862",
x"9E157803",
x"9CBD7783",
x"9B8476F5",
x"9A8E766E",
x"99FE760B",
x"99ED75E1",
x"9A677602",
x"9B6D7679",
x"9CF07743",
x"9ED67857",
x"A10179A3",
x"A34F7B12",
x"A5A17C91",
x"A7E17E09",
x"AA017F70",
x"ABF780BA",
x"ADC081E6",
x"AF6382F4",
x"B0E083E8",
x"B23984C6",
x"B36E858F",
x"B47E8643",
x"B56386DE",
x"B616875D",
x"B69C87B8",
x"B6F387EC",
x"B72087F3",
x"B73287CD",
x"B7358783",
x"B7368717",
x"B7438697",
x"B760860F",
x"B7928592",
x"B7D9852C",
x"B82C84ED",
x"B88584DD",
x"B8DB8502",
x"B9288560",
x"B96685EE",
x"B99286A4",
x"B9B5876E",
x"B9D1883C",
x"B9F188FB",
x"BA22899D",
x"BA6B8A14",
x"BAD78A5D",
x"BB688A7A",
x"BC1E8A71",
x"BCE88A4D",
x"BDB58A17",
x"BE5B89CF",
x"BEB08973",
x"BE7B88F0",
x"BD818832",
x"BB8B8718",
x"B86A8585",
x"B4048363",
x"AE5980A2",
x"A7857D4A",
x"9FC37971",
x"976C7540",
x"8EEA70F2",
x"86B56CC7",
x"7F3E68FF",
x"78E965D2",
x"74006366",
x"70A861CF",
x"6EE56108",
x"6E9760FE",
x"6F81618D",
x"71566287",
x"73C263C4",
x"7673651D",
x"79256679",
x"7BAA67C9",
x"7DE5690A",
x"7FD16A3F",
x"81746B70",
x"82E26CA1",
x"842F6DD5",
x"856F6F06",
x"86AA7029",
x"87E6712A",
x"891D71FB",
x"8A467289",
x"8B5372CD",
x"8C3972C1",
x"8CF1726E",
x"8D7771DF",
x"8DD3712D",
x"8E0B706C",
x"8E2F6FB3",
x"8E4D6F13",
x"8E716E9A",
x"8EA76E4E",
x"8EED6E2A",
x"8F456E27",
x"8FA56E3D",
x"90036E5B",
x"904D6E79",
x"90776E8D",
x"90716E92",
x"90326E85",
x"8FB26E66",
x"8EF36E3B",
x"8DFA6E06",
x"8CD06DCB",
x"8B896D8A",
x"8A346D48",
x"88E76D04",
x"87B86CC4",
x"86B76C86",
x"85F06C51",
x"856C6C28",
x"852B6C12",
x"85286C13",
x"855B6C2E",
x"85B46C66",
x"86276CBA",
x"86A76D23",
x"872A6D99",
x"87AC6E16",
x"882D6E8D",
x"88AF6EF9",
x"893C6F52",
x"89DC6F94",
x"8A946FC0",
x"8B676FD7",
x"8C556FDB",
x"8D536FD1",
x"8E556FC0",
x"8F496FAA",
x"901A6F92",
x"90B46F7A",
x"91066F64",
x"91016F4D",
x"90A26F34",
x"8FE76F1A",
x"8EDC6EFE",
x"8D8B6ED9",
x"8C0A6EAD",
x"8A706E75",
x"88D86E29",
x"87566DC7",
x"86076D4B",
x"84FB6CB4",
x"84456C02",
x"83EA6B3A",
x"83EF6A65",
x"844E6993",
x"84FB68D4",
x"85E66835",
x"86F967CB",
x"881B679D",
x"893967B5",
x"8A3E6813",
x"8B1B68B0",
x"8BCC6980",
x"8C4F6A75",
x"8CAC6B7D",
x"8CEC6C86",
x"8D206D80",
x"8D536E5E",
x"8D926F17",
x"8DE66FA6",
x"8E4D7008",
x"8EC3703B",
x"8F3E7044",
x"8FAC7021",
x"90016FD9",
x"902C6F70",
x"90246EEE",
x"8FE26E58",
x"8F666DBE",
x"8EB86D2B",
x"8DE56CB0",
x"8CF96C55",
x"8C046C26",
x"8B0E6C21",
x"8A1F6C45",
x"89326C80",
x"883F6CBE",
x"87356CE6",
x"86036CDE",
x"84976C8C",
x"82E46BE2",
x"80ED6ADB",
x"7EBA6983",
x"7C6567EF",
x"7A166645",
x"77FA64AD",
x"76466356",
x"752D626A",
x"74D5620D",
x"75546250",
x"76B2633B",
x"78DF64C4",
x"7BB766D1",
x"7F0B6941",
x"82A56BEB",
x"864C6EA6",
x"89CF714E",
x"8D0B73C8",
x"8FF075FF",
x"927B77EC",
x"94BE7993",
x"96D07AFC",
x"98D27C34",
x"9AE47D50",
x"9D1E7E5B",
x"9F8E7F65",
x"A2368078",
x"A50F819B",
x"A80A82CF",
x"AB0C8414",
x"AE018566",
x"B0DB86C5",
x"B38C882C",
x"B6148997",
x"B8778B04",
x"BABF8C6C",
x"BCFB8DC9",
x"BF368F13",
x"C175903C",
x"C3B79139",
x"C5F291FF",
x"C813927C",
x"CA0292AD",
x"CBA3928A",
x"CCDD921A",
x"CD9B9166",
x"CDD39081",
x"CD828F83",
x"CCB98E86",
x"CB898DA4",
x"CA138CF6",
x"C8788C87",
x"C6D48C60",
x"C5438C7A",
x"C3D78CC3",
x"C2958D25",
x"C17C8D81",
x"C0818DB8",
x"BF958DB1",
x"BEA88D58",
x"BDAF8CAA",
x"BCA58BAC",
x"BB8E8A71",
x"BA778917",
x"B97087BC",
x"B88B8683",
x"B7DD8587",
x"B76E84DD",
x"B740848D",
x"B74A8491",
x"B77B84DA",
x"B7B98552",
x"B7EB85DA",
x"B7FE865C",
x"B7E486C2",
x"B7A386FE",
x"B74A8714",
x"B6FB870A",
x"B6DD86F6",
x"B71986ED",
x"B7D7870A",
x"B92D8760",
x"BB2287FE",
x"BDA088E6",
x"C0828A0E",
x"C38B8B63",
x"C6728CCB",
x"C8F28E22",
x"CACB8F4C",
x"CBD3902F",
x"CBF790B9",
x"CB4190E2",
x"C9DA90B1",
x"C7FE9034",
x"C5F78F83",
x"C40C8EB9",
x"C27F8DF4",
x"C17E8D4B",
x"C11B8CD2",
x"C14A8C94",
x"C1F08C94",
x"C2D88CCF",
x"C3CC8D3E",
x"C4948DD3",
x"C5098E83",
x"C5188F41",
x"C4BC9001",
x"C40B90BC",
x"C3259165",
x"C23291F0",
x"C1509253",
x"C09B9280",
x"C016926A",
x"BFB99202",
x"BF6A913F",
x"BF06901B",
x"BE6A8E98",
x"BD7A8CC2",
x"BC268AAB",
x"BA75886C",
x"B87A8621",
x"B65683EA",
x"B43581E1",
x"B23B8016",
x"B0847E94",
x"AF187D4E",
x"ADE97C39",
x"ACD47B39",
x"ABA27A2D",
x"AA1578F9",
x"A7F3777F",
x"A50B75B1",
x"A142738B",
x"9C9B7116",
x"97366E6E",
x"91506BB2",
x"8B3C690E",
x"855366A8",
x"7FF764A3",
x"7B77631A",
x"7814621B",
x"75F261A5",
x"751661AE",
x"75696222",
x"76C262E9",
x"78E663E8",
x"7B91650A",
x"7E846641",
x"81886783",
x"847768CE",
x"87386A24",
x"89C56B8C",
x"8C256D0C",
x"8E696EA3",
x"90A47054",
x"92EA7217",
x"954C73E5",
x"97D275B3",
x"9A7B7777",
x"9D437928",
x"A01C7ABE",
x"A2F17C3C",
x"A5B27D9C",
x"A84C7EE1",
x"AAAC800F",
x"ACC98128",
x"AE9B822C",
x"B022831B",
x"B16183F6",
x"B26184BB",
x"B329856A",
x"B3C48604",
x"B43F868A",
x"B49E86FD",
x"B4E6875D",
x"B51487A9",
x"B52887DC",
x"B51987F0",
x"B4E187DD",
x"B47D879F",
x"B3E88732",
x"B3298698",
x"B24785D9",
x"B1548504",
x"B060842B",
x"AF7E8366",
x"AEC382C7",
x"AE388261",
x"ADE18239",
x"ADBC824C",
x"ADB9828F",
x"ADC382EB",
x"ADC38346",
x"AD9E8387",
x"AD3F8395",
x"AC9B8367",
x"ABAF82F7",
x"AA8A8251",
x"A940818A",
x"A7F580BD",
x"A6CF800C",
x"A5F37F92",
x"A5847F65",
x"A5977F94",
x"A638801C",
x"A76080F4",
x"A8FD8207",
x"AAEE8338",
x"AD11846A",
x"AF3C8585",
x"B1538676",
x"B33C872E",
x"B4ED87AC",
x"B66987FA",
x"B7BF8822",
x"B90A883C",
x"BA648859",
x"BBE8888E",
x"BDA988E9",
x"BFAF8974",
x"C1F28A31",
x"C4638B1E",
x"C6E28C32",
x"C9538D60",
x"CB928E9A",
x"CD868FCF",
x"CF1C90F3",
x"D04891F9",
x"D11092D6",
x"D1799386",
x"D1939403",
x"D16D944C",
x"D10F9462",
x"D0859448",
x"CFCE9400",
x"CEEC9390",
x"CDE09300",
x"CCA79253",
x"CB479191",
x"C9C790C1",
x"C8368FE5",
x"C6A08F01",
x"C5188E1B",
x"C3A68D35",
x"C2548C50",
x"C1258B73",
x"C0138AA4",
x"BF1B89EA",
x"BE308950",
x"BD4D88DF",
x"BC6E889F",
x"BB8F8894",
x"BAAF88BC",
x"B9CC8908",
x"B8DB8967",
x"B7D089B6",
x"B69189D0",
x"B4FD898D",
x"B2EE88C2",
x"B03F874F",
x"ACD3851C",
x"A8948229",
x"A3887E85",
x"9DC67A4D",
x"978175B9",
x"90FB7108",
x"8A8A6C7D",
x"84846862",
x"7F3F64EF",
x"7B026253",
x"77FD60AB",
x"764C5FFC",
x"75F06039",
x"76D26145",
x"78C462F6",
x"7B90651A",
x"7EF6677D",
x"82B569F0",
x"86936C4E",
x"8A5C6E76",
x"8DEA7058",
x"912271EE",
x"93F9733A",
x"96647448",
x"986E7527",
x"9A1F75E5",
x"9B847692",
x"9CAF7734",
x"9DAC77D4",
x"9E8A786E",
x"9F527901",
x"A0077981",
x"A0AF79EA",
x"A14A7A33",
x"A1D97A5E",
x"A25F7A6D",
x"A2DF7A6A",
x"A3637A64",
x"A3F77A6B",
x"A4A77A91",
x"A5827AE3",
x"A6947B67",
x"A7E47C1E",
x"A9717D01",
x"AB337DFF",
x"AD187F04",
x"AF0B7FFA",
x"B0ED80CA",
x"B2A18167",
x"B40B81C9",
x"B51481EE",
x"B5B281E1",
x"B5DE81B5",
x"B5A6817A",
x"B5188146",
x"B44E812C",
x"B36A8137",
x"B288816E",
x"B1C781CC",
x"B1408246",
x"B10082D0",
x"B1088354",
x"B15783C3",
x"B1D9840B",
x"B2748423",
x"B30A8404",
x"B37B83B1",
x"B3A8832C",
x"B3788287",
x"B2DE81CC",
x"B1D3810B",
x"B0618054",
x"AE9C7FB3",
x"ACA17F2F",
x"AA917ECD",
x"A8947E8A",
x"A6D07E60",
x"A5637E46",
x"A4667E33",
x"A3E67E20",
x"A3E47E07",
x"A4597DE5",
x"A5317DBF",
x"A6547D9B",
x"A7A67D82",
x"A90B7D7F",
x"AA677D9B",
x"ABA37DD7",
x"ACAD7E30",
x"AD777E9E",
x"ADFA7F0E",
x"AE307F6D",
x"AE187FA6",
x"ADB27FA3",
x"AD017F5A",
x"AC047EC1",
x"AAC27DDA",
x"A9407CAF",
x"A7877B51",
x"A5A279D7",
x"A39B7856",
x"A18476E1",
x"9F677589",
x"9D577455",
x"9B5F734B",
x"9988726A",
x"97D971AA",
x"9655710A",
x"94FA7085",
x"93C67016",
x"92B46FBD",
x"91BB6F76",
x"90D86F44",
x"90016F1E",
x"8F376F02",
x"8E706EE4",
x"8DAE6EBA",
x"8CEF6E78",
x"8C2F6E16",
x"8B706D8D",
x"8AB26CDF",
x"89F26C12",
x"892B6B30",
x"885C6A49",
x"877D6969",
x"8683689B",
x"855F67E3",
x"8401673B",
x"8258669A",
x"804F65EC",
x"7DD9651B",
x"7AEC6415",
x"778362CB",
x"73AA6134",
x"6F735F56",
x"6B005D43",
x"66765B15",
x"620658ED",
x"5DE256ED",
x"5A365536",
x"572953E3",
x"54D552FF",
x"5348528E",
x"52805287",
x"526C52D4",
x"52F2535E",
x"53F15409",
x"554554C0",
x"56CB556B",
x"58665604",
x"5A035687",
x"5B9656F8",
x"5D165761",
x"5E8957D0",
x"5FF2584C",
x"615658DD",
x"62BA5985",
x"641C5A3F",
x"65765B00",
x"66BF5BBC",
x"67EB5C63",
x"68E85CEA",
x"69AD5D48",
x"6A315D78",
x"6A705D7E",
x"6A705D64",
x"6A3B5D33",
x"69DF5CFD",
x"696D5CCF",
x"68F65CB6",
x"68875CB9",
x"682B5CDA",
x"67E65D17",
x"67B85D66",
x"679B5DBC",
x"678C5E0B",
x"67825E48",
x"677A5E66",
x"67735E62",
x"67725E39",
x"677C5DF3",
x"67995D9A",
x"67D25D3B",
x"682D5CE6",
x"68AB5CAE",
x"694B5C9C",
x"6A055CBC",
x"6ACB5D11",
x"6B905D97",
x"6C425E43",
x"6CD45F07",
x"6D385FD0",
x"6D6E6088",
x"6D6F611F",
x"6D456184",
x"6CFA61AE",
x"6C9D619A",
x"6C3F614B",
x"6BF260CE",
x"6BC46033",
x"6BC25F8D",
x"6BF25EF0",
x"6C585E6C",
x"6CF05E0D",
x"6DAF5DDA",
x"6E8C5DD5",
x"6F735DF6",
x"70565E35",
x"71235E84",
x"71C95ED7",
x"72425F27",
x"72895F69",
x"729E5F9D",
x"72895FC2",
x"72565FDD",
x"72145FF3",
x"71D2600A",
x"71A06025",
x"71866043",
x"718C6064",
x"71B16083",
x"71F06097",
x"723F609F",
x"72936095",
x"72DC607A",
x"7311604F",
x"732A601A",
x"73215FDF",
x"72FA5FA8",
x"72BB5F7A",
x"726C5F5A",
x"72185F49",
x"71CE5F46",
x"71965F4C",
x"71755F55",
x"71705F5A",
x"71875F5A",
x"71B55F52",
x"71F35F41",
x"72345F27",
x"72705F0A",
x"729A5EE9",
x"72AA5EC8",
x"72975EA5",
x"725C5E80",
x"71F75E55",
x"716C5E22",
x"70BA5DE6",
x"6FEC5D9C",
x"6F095D4B",
x"6E195CF1",
x"6D275C95",
x"6C3A5C3C",
x"6B535BE6",
x"6A775B95",
x"699E5B46",
x"68C25AF1",
x"67D85A8E",
x"66D25A12",
x"65A45975",
x"644758B3",
x"62B257CC",
x"60EB56C3",
x"5EF655A6",
x"5CE55481",
x"5ACA5367",
x"58BB5267",
x"56D2518F",
x"552350E7",
x"53C05072",
x"52B6502B",
x"520A5008",
x"51BE4FFF",
x"51C85005",
x"52215011",
x"52B9501C",
x"53825029",
x"546F503A",
x"5572505D",
x"56805099",
x"579050FB",
x"589D518C",
x"59A0524E",
x"5A97533F",
x"5B805454",
x"5C5B557E",
x"5D2A56AC",
x"5DF057C9",
x"5EB058BF",
x"5F6C597E",
x"602B59FD",
x"60EE5A36",
x"61B55A2C",
x"628359E7",
x"63575977",
x"642D58ED",
x"6503585D",
x"65D457D7",
x"6699576E",
x"674C572B",
x"67E95712",
x"68655725",
x"68BB575E",
x"68E357B5",
x"68DB581B",
x"689D5884",
x"682B58E3",
x"678D5933",
x"66CC5970",
x"65FA599B",
x"652B59BD",
x"647659E1",
x"63F25A14",
x"63B25A63",
x"63C85AD9",
x"643B5B7B",
x"650C5C49",
x"662E5D3B",
x"67915E41",
x"691E5F46",
x"6ABA6038",
x"6C4860FE",
x"6DB16187",
x"6EE361C8",
x"6FD461BC",
x"707F616F",
x"70E960EC",
x"7120604D",
x"71305FAE",
x"712D5F28",
x"71245ED5",
x"71245EC6",
x"71315F04",
x"714F5F8A",
x"717A604B",
x"71A86132",
x"71CF6222",
x"71E36300",
x"71DB63B1",
x"71B06423",
x"71616449",
x"70EF6427",
x"706563C5",
x"6FCB6338",
x"6F306297",
x"6EA061FC",
x"6E24617D",
x"6DC56129",
x"6D826107",
x"6D566114",
x"6D3B6141",
x"6D25617A",
x"6D0961A9",
x"6CDB61B7",
x"6C94618E",
x"6C336128",
x"6BBA6081",
x"6B315FA4",
x"6AA65EA4",
x"6A265D98",
x"69C15C9E",
x"69825BCF",
x"69725B3F",
x"69915AFD",
x"69DE5B08",
x"6A4E5B5D",
x"6AD25BE9",
x"6B5F5C95",
x"6BE25D4B",
x"6C4E5DF0",
x"6C9A5E6E",
x"6CC15EB9",
x"6CC25EC9",
x"6CA45E9E",
x"6C6D5E41",
x"6C275DBF",
x"6BDE5D28",
x"6B975C90",
x"6B5C5C02",
x"6B305B90",
x"6B105B3C",
x"6AFA5B0D",
x"6AE55AFD",
x"6AC75B08",
x"6A945B24",
x"6A415B42",
x"69C55B5A",
x"69175B5F",
x"68345B47",
x"671B5B10",
x"65D55AB5",
x"646C5A39",
x"62F359A2",
x"618258FA",
x"602E584A",
x"5F1357A2",
x"5E47570E",
x"5DDB569B",
x"5DDC5653",
x"5E4D5640",
x"5F295667",
x"606556C6",
x"61EF575C",
x"63B4581E",
x"659E5904",
x"679A5A01",
x"699C5B08",
x"6B975C10",
x"6D895D0B",
x"6F725DF8",
x"71565ED2",
x"733E5F9B",
x"752B605A",
x"7727611A",
x"793161E3",
x"7B4E62C5",
x"7D7663C6",
x"7FA864F2",
x"81DB6648",
x"840667C5",
x"861D695F",
x"88176B07",
x"89E66CA8",
x"8B806E2D",
x"8CE06F7F",
x"8DFE708A",
x"8EDA7143",
x"8F76719F",
x"8FD971A1",
x"90107155",
x"902470CA",
x"90247014",
x"901B6F4F",
x"90136E92",
x"90116DF0",
x"90156D7C",
x"901F6D3B",
x"902B6D34",
x"90326D62",
x"90326DBE",
x"902E6E3E",
x"90286ED5",
x"902B6F79",
x"90417021",
x"907770C5",
x"90D9715F",
x"916F71EF",
x"92397274",
x"933672EC",
x"945A735A",
x"959573BE",
x"96D3741A",
x"97FE746F",
x"990474BD",
x"99D27503",
x"9A5D7546",
x"9A9F757F",
x"9A9575B0",
x"9A4675D5",
x"99B875EE",
x"98F975F4",
x"981775E5",
x"972175BE",
x"962B7581",
x"9545752C",
x"948074C7",
x"93EC7457",
x"939273E6",
x"937B737F",
x"93A8732D",
x"941272F9",
x"94AC72E8",
x"956472FE",
x"961F7336",
x"96C3738B",
x"973873EE",
x"976A7454",
x"974B74AD",
x"96D974EA",
x"961C74FF",
x"952574E5",
x"940A749A",
x"92E67421",
x"91D37382",
x"90E472C4",
x"902B71F6",
x"8FAB7127",
x"8F637062",
x"8F466FB4",
x"8F4B6F29",
x"8F606EC4",
x"8F7A6E8D",
x"8F906E89",
x"8F9E6EB4",
x"8FA96F0D",
x"8FB96F90",
x"8FD97035",
x"901170F6",
x"906E71C7",
x"90F4729F",
x"91A77374",
x"9283743E",
x"938174F9",
x"949B75A2",
x"95BF7639",
x"96E376BE",
x"97F77739",
x"98ED77AC",
x"99B9781B",
x"9A527889",
x"9AB178F4",
x"9ACF7956",
x"9AAE79A8",
x"9A4D79DB",
x"99AF79E3",
x"98D379B0",
x"97B97933",
x"965A7860",
x"94AE772C",
x"92A77593",
x"90397397",
x"8D5B7143",
x"8A076EA1",
x"86436BCE",
x"822568E2",
x"7DCF65FF",
x"79706348",
x"754760DD",
x"718D5EE0",
x"6E845D69",
x"6C5E5C84",
x"6B3A5C3B",
x"6B245C87",
x"6C135D5A",
x"6DE65E9F",
x"706B6038",
x"73686207",
x"76A063ED",
x"79DC65CF",
x"7CF36799",
x"7FC8693A",
x"824F6AAA",
x"848A6BE9",
x"86866CFA",
x"88536DE6",
x"8A066EB4",
x"8BA86F6F",
x"8D43701D",
x"8ED970C8",
x"90647172",
x"91DF721A",
x"933F72C1",
x"94817364",
x"95A573FE",
x"96AC7489",
x"979D7503",
x"98807568",
x"995D75B9",
x"9A3875F1",
x"9B107616",
x"9BE37627",
x"9CA47629",
x"9D48761D",
x"9DBF7605",
x"9DFB75E4",
x"9DF375BC",
x"9DA2758C",
x"9D0A7558",
x"9C317523",
x"9B2674F1",
x"99FB74C6",
x"98C274A7",
x"978E749C",
x"967074A6",
x"957474C4",
x"94A174F6",
x"93F77536",
x"93767576",
x"931875AF",
x"92D975D2",
x"92B475D8",
x"92A475BA",
x"92A87578",
x"92C57516",
x"92FB74A3",
x"9352742D",
x"93CB73C6",
x"9463737C",
x"9518735E",
x"95E27372",
x"96B173B9",
x"97777429",
x"982274B4",
x"98A2754A",
x"98EE75D5",
x"98FE7644",
x"98D67689",
x"9881769F",
x"98117683",
x"979B763E",
x"973875DE",
x"96FD756F",
x"96FB7506",
x"973C74AF",
x"97BF7475",
x"9879745C",
x"99557462",
x"9A397480",
x"9B0874AA",
x"9BA674D4",
x"9BFD74EF",
x"9BFD74F5",
x"9BA574DE",
x"9AFB74AD",
x"9A127464",
x"9903740F",
x"97E673B7",
x"96DA736B",
x"95F87333",
x"954F7317",
x"94E6731C",
x"94C17343",
x"94D27386",
x"951173E2",
x"956A744B",
x"95CF74BA",
x"96317523",
x"9684757C",
x"96C575BC",
x"96EE75DA",
x"970175D0",
x"96FB7596",
x"96E0752D",
x"96A97492",
x"965573CA",
x"95DD72DC",
x"953F71D7",
x"947670CA",
x"93886FCA",
x"927E6EE9",
x"91666E3D",
x"90566DD2",
x"8F606DB3",
x"8E986DDC",
x"8E0A6E41",
x"8DB56ECD",
x"8D8B6F5F",
x"8D716FD2",
x"8D3C7000",
x"8CBB6FC5",
x"8BBE6F08",
x"8A176DB7",
x"87AA6BD4",
x"8471696F",
x"807E66AA",
x"7C0163B5",
x"773C60C3",
x"72845E12",
x"6E345BD5",
x"6AA15A36",
x"68135955",
x"66B8593C",
x"66A359E6",
x"67C75B39",
x"69FD5D14",
x"6D095F49",
x"70A461A9",
x"7487640A",
x"78736645",
x"7C386844",
x"7FBB69F6",
x"82F46B5C",
x"85EA6C7C",
x"88B16D68",
x"8B606E2E",
x"8E0D6EE4",
x"90C26F99",
x"9380705A",
x"963C712D",
x"98DF7215",
x"9B4F730F",
x"9D6E7413",
x"9F27751D",
x"A06A7620",
x"A1367713",
x"A19777EF",
x"A19E78AC",
x"A16B7944",
x"A12279B9",
x"A0E37A0C",
x"A0CC7A43",
x"A0F47A68",
x"A16A7A89",
x"A22E7AB2",
x"A3367AED",
x"A46D7B43",
x"A5B67BB4",
x"A6EA7C3D",
x"A7E07CCE",
x"A86D7D56",
x"A86A7DB9",
x"A7B87DE0",
x"A6427DB0",
x"A4057D1B",
x"A10F7C18",
x"9D7E7AAD",
x"998478EB",
x"955C76EB",
x"914874D2",
x"8D8A72C5",
x"8A5D70EB",
x"87EA6F5E",
x"86486E34",
x"85766D75",
x"85606D1D",
x"85DF6D1D",
x"86BC6D5C",
x"87C26DC1",
x"88B86E31",
x"89736E96",
x"89D66EE1",
x"89D56F0C",
x"89746F17",
x"88CB6F0D",
x"87F76EFC",
x"871E6EEF",
x"86606EF5",
x"85D66F13",
x"858E6F4D",
x"85876F9C",
x"85B26FF8",
x"85F6704F",
x"86347096",
x"864970BA",
x"862170B3",
x"85AF707A",
x"84FA7017",
x"841A6F93",
x"83376F02",
x"82896E7C",
x"824C6E1C",
x"82B86DFD",
x"83F76E35",
x"86216ED5",
x"892F6FE2",
x"8D047158",
x"91647329",
x"9601753B",
x"9A847771",
x"9E9479A6",
x"A1E67BB7",
x"A4467D87",
x"A5987EFA",
x"A5E37FFE",
x"A545808E",
x"A3F480A9",
x"A236805B",
x"A0527FB2",
x"9E877EC4",
x"9D087DA5",
x"9BF37C6A",
x"9B527B25",
x"9B1879E4",
x"9B2978B4",
x"9B64779B",
x"9B9B7699",
x"9BAC75AD",
x"9B7774D5",
x"9AEB740C",
x"9A04734E",
x"98C97297",
x"974D71E8",
x"95A57140",
x"93ED709D",
x"92387003",
x"90946F70",
x"8F066EE4",
x"8D866E57",
x"8BFE6DC2",
x"8A586D1A",
x"886F6C51",
x"86276B59",
x"83666A28",
x"802068B4",
x"7C5866FA",
x"78246503",
x"73AA62D9",
x"6F216093",
x"6AC85E4C",
x"66E25C22",
x"63AE5A36",
x"615F58A4",
x"60165782",
x"5FE256E1",
x"60BA56C6",
x"6282572E",
x"650A580A",
x"681A594A",
x"6B785AD6",
x"6EE85C95",
x"72385E70",
x"75476053",
x"7800622F",
x"7A5F63FC",
x"7C7365B2",
x"7E536755",
x"801E68E6",
x"81F96A70",
x"84016BF6",
x"86506D83",
x"88F66F19",
x"8BF670BB",
x"8F48726C",
x"92D97426",
x"968E75E2",
x"9A4A7798",
x"9DEA793A",
x"A14F7ABE",
x"A4607C15",
x"A70A7D32",
x"A93F7E0B",
x"AAFB7E9E",
x"AC3F7EE8",
x"AD117EEE",
x"AD787EBD",
x"AD857E63",
x"AD437DEF",
x"ACBF7D77",
x"AC047D08",
x"AB217CB2",
x"AA227C77",
x"A9167C5B",
x"A80D7C59",
x"A7117C63",
x"A6307C6E",
x"A5767C71",
x"A4E47C5E",
x"A4817C32",
x"A44A7BED",
x"A43B7B95",
x"A4467B36",
x"A4637ADD",
x"A4817A96",
x"A4957A6F",
x"A4927A6F",
x"A46E7A95",
x"A4247ADD",
x"A3AE7B3A",
x"A3117BA0",
x"A2537BFC",
x"A17D7C41",
x"A09E7C63",
x"9FC67C56",
x"9F077C1C",
x"9E737BB9",
x"9E1B7B33",
x"9E087A9C",
x"9E4579FF",
x"9ED0796F",
x"9FA478F9",
x"A0B478A9",
x"A1EE7888",
x"A33D789B",
x"A48E78DE",
x"A5C97951",
x"A6E079EB",
x"A7C67AA0",
x"A8787B64",
x"A8F57C29",
x"A9467CE5",
x"A9717D8C",
x"A9847E16",
x"A9887E81",
x"A98A7ECC",
x"A98C7EF7",
x"A9987F0A",
x"A9AB7F0A",
x"A9C57EFE",
x"A9E07EED",
x"A9F67ED1",
x"AA007EB0",
x"A9F07E81",
x"A9BD7E3D",
x"A95D7DDB",
x"A8C37D54",
x"A7EA7CA2",
x"A6CC7BC3",
x"A56D7ABA",
x"A3D67993",
x"A217785B",
x"A0457726",
x"9E787606",
x"9CC9750F",
x"9B4B744D",
x"9A0A73C8",
x"990D7383",
x"984C7375",
x"97BC7395",
x"974673D0",
x"96D77417",
x"9657745B",
x"95B8748C",
x"94F174A3",
x"9406749C",
x"92F77474",
x"91D3742C",
x"90A273C3",
x"8F6C7339",
x"8E2F7289",
x"8CE971AD",
x"8B8A70A1",
x"8A066F5E",
x"88536DE5",
x"866C6C41",
x"845C6A80",
x"823768BE",
x"8020671D",
x"7E4465C1",
x"7CD564CC",
x"7C01645D",
x"7BF06487",
x"7CB5654E",
x"7E5866A7",
x"80C86879",
x"83E56AA4",
x"87816D00",
x"8B706F66",
x"8F7E71B9",
x"938473E1",
x"976975D2",
x"9B1E7793",
x"9EAB7930",
x"A21B7ABC",
x"A5887C4D",
x"A90C7DF4",
x"ACBF7FBD",
x"B0AC81AD",
x"B4DC83BF",
x"B94285E4",
x"BDC68808",
x"C24A8A14",
x"C6A28BF4",
x"CAA58D95",
x"CE2C8EED",
x"D1188FF9",
x"D35A90BB",
x"D4EF9141",
x"D5EE919B",
x"D67491E0",
x"D6B39228",
x"D6DE9289",
x"D72A9311",
x"D7C893D2",
x"D8D894CC",
x"DA6595FD",
x"DC6C9759",
x"DED098CB",
x"E1679A3B",
x"E3F99B90",
x"E6529CB0",
x"E83D9D88",
x"E9909E0C",
x"EA379E38",
x"EA2D9E16",
x"E9809DB4",
x"E84E9D2C",
x"E6BB9C92",
x"E4F69C00",
x"E3269B8A",
x"E16E9B3A",
x"DFE79B15",
x"DE9F9B13",
x"DD9A9B27",
x"DCD59B41",
x"DC449B48",
x"DBD79B2D",
x"DB7E9ADB",
x"DB279A4C",
x"DAC3997B",
x"DA40986B",
x"D9959729",
x"D8B695C5",
x"D79D9455",
x"D64E92F2",
x"D4D091B4",
x"D33390B2",
x"D18C9003",
x"CFF78FB1",
x"CE928FC6",
x"CD78903E",
x"CCBF910A",
x"CC6F921A",
x"CC88934F",
x"CCF7948A",
x"CDA295AD",
x"CE619699",
x"CF0E973A",
x"CF829782",
x"CFA2976E",
x"CF5D9707",
x"CEB0965E",
x"CDAC9587",
x"CC6A9499",
x"CB0993AA",
x"C9AF92C9",
x"C87791FD",
x"C7719148",
x"C6A690A2",
x"C60C9000",
x"C5908F51",
x"C51B8E8A",
x"C48C8DA2",
x"C3D08C97",
x"C2D78B6C",
x"C1A38A2B",
x"C03F88E9",
x"BEC787B6",
x"BD6086A9",
x"BC2D85D3",
x"BB578543",
x"BAFB8500",
x"BB2B850D",
x"BBE48564",
x"BD1E85FD",
x"BEB686C9",
x"C08B87BB",
x"C26E88C3",
x"C43789D6",
x"C5C68AEA",
x"C7058BF6",
x"C7F28CF9",
x"C8968DF1",
x"C90B8EE0",
x"C96F8FC5",
x"C9E0909D",
x"CA6F9160",
x"CB259203",
x"CBEB9270",
x"CC96928E",
x"CCE49244",
x"CC7E916D",
x"CB0E8FF3",
x"C83F8DBE",
x"C3D18AC3",
x"BDA68708",
x"B5C982A1",
x"AC747DB2",
x"A208786B",
x"970E730C",
x"8C206DD4",
x"81E26904",
x"78E764D6",
x"71AB6177",
x"6C7C5F00",
x"697B5D7A",
x"68935CD9",
x"69875D02",
x"6BFA5DD2",
x"6F7A5F18",
x"739060AB",
x"77CF6260",
x"7BDE641B",
x"7F8365C8",
x"82A1675F",
x"853868E3",
x"875F6A61",
x"893E6BE3",
x"8AFD6D7C",
x"8CC86F30",
x"8EB87100",
x"90E072E8",
x"933B74D7",
x"95B976B9",
x"98407877",
x"9AAC79FB",
x"9CDC7B34",
x"9EB27C18",
x"A01B7CA3",
x"A1117CDE",
x"A1977CD7",
x"A1BF7CA2",
x"A1A47C53",
x"A15F7BFE",
x"A1117BB6",
x"A0D47B85",
x"A0BB7B6E",
x"A0CF7B74",
x"A1127B92",
x"A1807BBF",
x"A2087BF4",
x"A29E7C2C",
x"A32C7C60",
x"A3A57C8F",
x"A3F87CB9",
x"A41E7CDD",
x"A40F7CF7",
x"A3CF7D06",
x"A35D7D06",
x"A2C37CF2",
x"A20D7CC3",
x"A1467C74",
x"A0817C05",
x"9FCD7B78",
x"9F387AD4",
x"9ECC7A23",
x"9E8F7972",
x"9E8478CB",
x"9EA27839",
x"9EDA77BE",
x"9F18775D",
x"9F42770C",
x"9F3F76C3",
x"9EF87674",
x"9E5D7612",
x"9D6A7593",
x"9C2274F8",
x"9A977446",
x"98E37386",
x"972972D0",
x"958E7237",
x"943671D5",
x"933F71BA",
x"92BC71F0",
x"92B67279",
x"932B734B",
x"94087451",
x"9535756F",
x"96947686",
x"9801777B",
x"995F7833",
x"9A91789C",
x"9B8478B3",
x"9C2F787B",
x"9C907802",
x"9CA9775E",
x"9C8A76A7",
x"9C3D75F9",
x"9BD67565",
x"9B6174FE",
x"9AEA74C7",
x"9A7674C3",
x"9A0574E7",
x"999A7525",
x"9929756B",
x"98AF75AA",
x"982575D0",
x"978775D1",
x"96D375A7",
x"96107554",
x"954374DA",
x"94797446",
x"93BB73A5",
x"93147306",
x"928B7275",
x"922271FE",
x"91D871A6",
x"91A1716B",
x"9176714B",
x"9149713A",
x"9111712D",
x"90C57117",
x"906470EE",
x"8FF270AA",
x"8F737048",
x"8EF06FCA",
x"8E716F34",
x"8DFD6E8F",
x"8D906DDF",
x"8D1D6D2A",
x"8C946C70",
x"8BD96BB0",
x"8ACE6ADE",
x"895669F5",
x"875D68E9",
x"84D567B5",
x"81C26658",
x"7E3B64D6",
x"7A63633B",
x"7670619A",
x"72A0600A",
x"6F2E5EA5",
x"6C595D81",
x"6A525CB5",
x"69385C4F",
x"69195C56",
x"69EB5CC8",
x"6B965D9C",
x"6DF05EC3",
x"70C86028",
x"73E861B4",
x"771D6350",
x"7A3B64E6",
x"7D236663",
x"7FBE67BA",
x"820468E3",
x"83F969DC",
x"85A26AA7",
x"87106B4C",
x"88536BD5",
x"89796C4D",
x"8A916CBF",
x"8BA76D3A",
x"8CBF6DC1",
x"8DDD6E5B",
x"8F066F06",
x"90356FC3",
x"91697088",
x"929D7151",
x"93C97217",
x"94E772D2",
x"95EE737E",
x"96D57416",
x"9790749A",
x"98177509",
x"98647562",
x"987475A7",
x"984975D7",
x"97E975F1",
x"975C75F4",
x"96B275DE",
x"95FA75B1",
x"9542756C",
x"94987513",
x"940874AC",
x"939A743D",
x"934D73D1",
x"93257375",
x"931F7333",
x"93387316",
x"936F7327",
x"93C8736E",
x"944873EB",
x"94F6749D",
x"95DF757C",
x"9708767F",
x"987B7795",
x"9A3478AC",
x"9C2C79AF",
x"9E507A8E",
x"A0887B36",
x"A2B37B9F",
x"A4AC7BC1",
x"A6507BA0",
x"A7817B46",
x"A8267AC0",
x"A8367A23",
x"A7AF7983",
x"A69E78F2",
x"A5187881",
x"A33B7834",
x"A126780C",
x"9EFD7803",
x"9CD9780B",
x"9AD67813",
x"9907780F",
x"977677EF",
x"962C77B0",
x"952E7751",
x"947776D8",
x"94077652",
x"93D775CB",
x"93E17554",
x"941B74F4",
x"947974B1",
x"94EC748D",
x"95647485",
x"95CF748D",
x"961A749D",
x"963874AA",
x"961F74AF",
x"95C874A5",
x"9536748D",
x"94717468",
x"938B743A",
x"92957408",
x"91A773D1",
x"90D67397",
x"9037735B",
x"8FD9731C",
x"8FC572DB",
x"8FFC7299",
x"9076725B",
x"9125722A",
x"91F6720C",
x"92D2720A",
x"939E722B",
x"9445726C",
x"94B172CB",
x"94D3733B",
x"94A873AF",
x"942E7410",
x"936F7450",
x"927B745C",
x"916C742D",
x"905273BE",
x"8F487319",
x"8E597245",
x"8D907157",
x"8CE9705C",
x"8C586F66",
x"8BC56E80",
x"8B136DAD",
x"8A246CE8",
x"88D96C27",
x"871B6B5E",
x"84E26A7A",
x"822E6975",
x"7F176846",
x"7BBF66F2",
x"78566586",
x"75146415",
x"723562BE",
x"6FED619D",
x"6E6860CF",
x"6DC1606C",
x"6E046083",
x"6F286117",
x"71136222",
x"739E6391",
x"769B6549",
x"79D8672D",
x"7D27691B",
x"80636AFA",
x"83746CB5",
x"86526E44",
x"88FE6FA1",
x"8B8970D8",
x"8E0471F5",
x"908B7308",
x"932F7423",
x"96007552",
x"990376A0",
x"9C2F780C",
x"9F787990",
x"A2C27B25",
x"A5F07CB6",
x"A8E17E36",
x"AB777F91",
x"AD9480B6",
x"AF288198",
x"B026822B",
x"B08C8268",
x"B0608253",
x"AFB081ED",
x"AE948142",
x"AD258060",
x"AB847F5A",
x"A9CC7E49",
x"A8217D3D",
x"A6997C50",
x"A54D7B92",
x"A4497B0E",
x"A3907AC7",
x"A31E7ABC",
x"A2E67AE1",
x"A2D77B28",
x"A2DF7B79",
x"A2E67BC6",
x"A2E17BFC",
x"A2CA7C12",
x"A29F7C06",
x"A26A7BE0",
x"A23C7BA8",
x"A2267B74",
x"A2387B53",
x"A27D7B58",
x"A2F77B8F",
x"A39C7BF7",
x"A4597C8B",
x"A50E7D3C",
x"A59E7DEF",
x"A5E67E8E",
x"A5CF7EFC",
x"A54C7F26",
x"A4617F01",
x"A3267E8C",
x"A1BF7DD1",
x"A05F7CEB",
x"9F3F7BF8",
x"9E927B1E",
x"9E877A81",
x"9F387A40",
x"A0A87A6E",
x"A2C67B13",
x"A56A7C28",
x"A85C7D94",
x"AB567F36",
x"AE1580EB",
x"B064828B",
x"B21683F4",
x"B318850B",
x"B36D85C6",
x"B3308622",
x"B28B862C",
x"B1AC85F4",
x"B0C58591",
x"AFFB8517",
x"AF668499",
x"AF0A8421",
x"AEDA83B2",
x"AEBD834C",
x"AE9182E8",
x"AE368282",
x"AD9B8219",
x"ACB881AF",
x"AB98814A",
x"AA5A80F7",
x"A92580C0",
x"A82580AD",
x"A78180C5",
x"A7538100",
x"A7A58153",
x"A86981AC",
x"A98081F4",
x"AAB98211",
x"ABE081F0",
x"ACC08185",
x"AD2E80CF",
x"AD127FD1",
x"AC677EA3",
x"AB3C7D5A",
x"A9B37C12",
x"A7FA7AE8",
x"A63F79F2",
x"A4AF793C",
x"A36778C8",
x"A273788F",
x"A1C9787C",
x"A1487875",
x"A0C07856",
x"9FF377FB",
x"9E9F7746",
x"9C877617",
x"997A7462",
x"955D721F",
x"90316F57",
x"8A116C21",
x"833768A3",
x"7BF6650A",
x"74AF618A",
x"6DCF5E57",
x"67BF5BA4",
x"62DB5994",
x"5F665842",
x"5D8957B5",
x"5D4857E6",
x"5E8958BC",
x"61175A18",
x"64A45BCF",
x"68DB5DB9",
x"6D655FB1",
x"71F36197",
x"764A6356",
x"7A3D64E6",
x"7DBB6642",
x"80C5676F",
x"83686876",
x"85BB695F",
x"87D86A32",
x"89D86AF7",
x"8BC96BB7",
x"8DB86C75",
x"8FA76D3A",
x"91976E10",
x"93846F02",
x"956C701D",
x"974F716C",
x"993272F9",
x"9B1874C6",
x"9D0776CB",
x"9F0378FC",
x"A1077B41",
x"A3117D7E",
x"A5157F8F",
x"A7038159",
x"A8CA82BD",
x"AA5C83AF",
x"ABAD8425",
x"ACB88426",
x"AD7B83C3",
x"ADFF8315",
x"AE528237",
x"AE7D814C",
x"AE8C8068",
x"AE8C7FA2",
x"AE7F7F05",
x"AE677E92",
x"AE427E43",
x"AE077E0E",
x"ADB27DE5",
x"AD407DBC",
x"ACB37D8B",
x"AC0C7D4D",
x"AB577D05",
x"AAA17CBA",
x"A9F67C75",
x"A9647C41",
x"A8F47C26",
x"A8A87C29",
x"A87B7C47",
x"A8637C7A",
x"A8507CB4",
x"A82F7CE7",
x"A7ED7D01",
x"A77A7CF2",
x"A6CF7CB2",
x"A5ED7C3F",
x"A4E37BA2",
x"A3C57AEA",
x"A2B37A30",
x"A1D27992",
x"A140792C",
x"A11B7912",
x"A16E7957",
x"A23D79F9",
x"A3777AF2",
x"A4FB7C25",
x"A6A57D72",
x"A8427EB5",
x"A9A67FC2",
x"AAAE807E",
x"AB4080D4",
x"AB5980BF",
x"AB028046",
x"AA577F82",
x"A97E7E96",
x"A89F7DA5",
x"A7DF7CD0",
x"A7597C36",
x"A71B7BE5",
x"A7247BE5",
x"A7637C2C",
x"A7BC7CA8",
x"A80F7D40",
x"A83F7DDE",
x"A8337E6E",
x"A7E37EE0",
x"A7527F2F",
x"A6947F60",
x"A5CC7F7C",
x"A51F7F91",
x"A4B87FA9",
x"A4B87FD3",
x"A5398015",
x"A6458071",
x"A7D780E3",
x"A9DA8166",
x"AC2C81F1",
x"AEA2827D",
x"B1158301",
x"B35E837E",
x"B56183F4",
x"B70A8464",
x"B85484D6",
x"B949854C",
x"B9F485CA",
x"BA68864F",
x"BAB086D3",
x"BAD4874D",
x"BACA87A8",
x"BA7B87D0",
x"B9C387A9",
x"B8758717",
x"B65E8600",
x"B34F844D",
x"AF2881F4",
x"A9DA7EF4",
x"A3717B54",
x"9C157731",
x"940B72B3",
x"8BB16E09",
x"836F696F",
x"7BB76523",
x"74F4615C",
x"6F835E4C",
x"6BA75C1A",
x"69825AD7",
x"691A5A8A",
x"6A515B1F",
x"6CF25C7A",
x"70B15E6E",
x"753C60CF",
x"7A3D6368",
x"7F65660D",
x"84736899",
x"89396AF5",
x"8D9A6D12",
x"918B6EF0",
x"9510709A",
x"9833721C",
x"9B087389",
x"9DA174F1",
x"A00B765B",
x"A24D77CB",
x"A469793D",
x"A6567AA3",
x"A80B7BEB",
x"A97E7D06",
x"AAA17DE5",
x"AB707E7C",
x"ABEA7ECF",
x"AC187EE4",
x"AC087ECD",
x"ABD07EA2",
x"AB877E7B",
x"AB457E70",
x"AB1F7E92",
x"AB237EEA",
x"AB597F75",
x"ABBC802B",
x"AC4280F4",
x"ACD681BD",
x"AD64826D",
x"ADD682ED",
x"AE188332",
x"AE198335",
x"ADD482F7",
x"AD4C8284",
x"AC8881E8",
x"AB978137",
x"AA8C8082",
x"A9807FD7",
x"A8817F40",
x"A7A17EC7",
x"A6ED7E6D",
x"A66B7E36",
x"A61C7E22",
x"A6007E30",
x"A60E7E5D",
x"A63F7EA5",
x"A6857F01",
x"A6D77F6A",
x"A7287FD3",
x"A769802F",
x"A7918072",
x"A797808F",
x"A7758080",
x"A72E8042",
x"A6C37FDA",
x"A6457F56",
x"A5BF7EC7",
x"A5467E3D",
x"A4ED7DCA",
x"A4C27D7B",
x"A4CF7D56",
x"A5187D56",
x"A5917D71",
x"A62C7D98",
x"A6CD7DB5",
x"A7567DB6",
x"A7AB7D8E",
x"A7AF7D35",
x"A7507CAF",
x"A68A7C02",
x"A5627B41",
x"A3EA7A7E",
x"A23D79CA",
x"A0807933",
x"9ED478C3",
x"9D597879",
x"9C267853",
x"9B467844",
x"9AB87841",
x"9A70783C",
x"9A5A7827",
x"9A5D77FF",
x"9A6377C0",
x"9A57776A",
x"9A347703",
x"99F97695",
x"99B17626",
x"997075C1",
x"994D7571",
x"9960753B",
x"99B97527",
x"9A637536",
x"9B567568",
x"9C8475BC",
x"9DD57627",
x"9F2576A6",
x"A056772C",
x"A14A77AD",
x"A1EE7820",
x"A23F7882",
x"A23F78CB",
x"A2057903",
x"A1AC792D",
x"A1507954",
x"A10A7982",
x"A0E979BD",
x"A0EA7A08",
x"A0FA7A5D",
x"A0F57AAC",
x"A0AB7AE0",
x"9FE67ADA",
x"9E6E7A7B",
x"9C2279A9",
x"98E97853",
x"94CD7671",
x"8FEE7410",
x"8A8A714A",
x"84F16E4B",
x"7F836B45",
x"7A9D6875",
x"769A660D",
x"73BB643C",
x"7230631F",
x"720262C4",
x"7325631F",
x"756F641D",
x"78A16595",
x"7C73675F",
x"8098694E",
x"84C86B3A",
x"88C36D06",
x"8C5D6E9D",
x"8F796FFE",
x"92097127",
x"940D7229",
x"95957310",
x"96B273EB",
x"977D74C6",
x"980D75A2",
x"98797681",
x"98D07758",
x"99277820",
x"998478CE",
x"99F1795A",
x"9A7379BD",
x"9B0B79F8",
x"9BBB7A12",
x"9C7D7A15",
x"9D4D7A0B",
x"9E2279FF",
x"9EF179FB",
x"9FAF7A03",
x"A04C7A19",
x"A0B97A36",
x"A0EE7A51",
x"A0E07A61",
x"A08D7A5D",
x"9FF67A3C",
x"9F2579FB",
x"9E29799D",
x"9D187925",
x"9C06789D",
x"9B07780D",
x"9A317782",
x"99917702",
x"992E7690",
x"99047630",
x"990D75E1",
x"9936759F",
x"996D7567",
x"999B7539",
x"99AB7510",
x"998E74F2",
x"993C74DC",
x"98B174D4",
x"97F174D7",
x"970874E2",
x"960374F2",
x"94EC74FB",
x"93D274F4",
x"92B974D1",
x"91A97486",
x"90A1740D",
x"8F9A7366",
x"8E927293",
x"8D86719F",
x"8C717099",
x"8B5C6F90",
x"8A4C6E99",
x"894C6DC1",
x"886A6D16",
x"87B56C9C",
x"87376C57",
x"86F46C3F",
x"86F36C4E",
x"872A6C78",
x"878E6CB0",
x"88136CEC",
x"88A56D23",
x"89386D4B",
x"89BB6D63",
x"8A276D66",
x"8A746D54",
x"8AA46D2D",
x"8AB66CF3",
x"8AB26CA8",
x"8A9A6C52",
x"8A736BF5",
x"8A426B96",
x"8A096B3B",
x"89CC6AEF",
x"898E6AB5",
x"89566A99",
x"89286A9C",
x"890D6AC2",
x"890B6B0D",
x"89296B79",
x"896A6C02",
x"89CF6CA3",
x"8A506D4F",
x"8AE76E02",
x"8B836EAE",
x"8C156F48",
x"8C8E6FC5",
x"8CDF701C",
x"8CFA7041",
x"8CDF702D",
x"8C8D6FDE",
x"8C0D6F52",
x"8B6D6E92",
x"8ABE6DA6",
x"8A106C9E",
x"89726B8F",
x"88EC6A89",
x"887C699E",
x"881568D9",
x"87A5683C",
x"870D67C2",
x"8628675C",
x"84D266F3",
x"82ED666D",
x"806665B4",
x"7D3A64B5",
x"79776368",
x"754861D3",
x"70E1600B",
x"6C8D5E31",
x"68975C70",
x"654F5AF3",
x"62F659E6",
x"61BA5969",
x"61B4598F",
x"62DE5A5C",
x"651A5BC0",
x"68375D9F",
x"6BF25FD3",
x"70056231",
x"742E648D",
x"783466C6",
x"7BEF68C2",
x"7F486A76",
x"823B6BDF",
x"84CF6D09",
x"87186E02",
x"892F6EDC",
x"8B2C6FAD",
x"8D257083",
x"8F277168",
x"9139725F",
x"9362736A",
x"959A747E",
x"97DC7595",
x"9A1B76A3",
x"9C4C779D",
x"9E5D787C",
x"A0427936",
x"A1E979C4",
x"A3497A26",
x"A4567A5B",
x"A50D7A67",
x"A5717A4E",
x"A58E7A1C",
x"A57379DA",
x"A5337995",
x"A4E97957",
x"A4A9792D",
x"A485791C",
x"A488792A",
x"A4B67957",
x"A508799D",
x"A57679F4",
x"A5EE7A51",
x"A6637AAD",
x"A6C97AFE",
x"A71B7B40",
x"A7567B72",
x"A7817B99",
x"A7A57BBC",
x"A7CC7BE3",
x"A8017C16",
x"A8467C5D",
x"A89E7CB7",
x"A9017D26",
x"A9677D9F",
x"A9C57E19",
x"AA0F7E85",
x"AA3D7ED9",
x"AA4C7F07",
x"AA3B7F0E",
x"AA0C7EF0",
x"A9CA7EAC",
x"A97A7E51",
x"A9247DED",
x"A8CD7D8E",
x"A87D7D43",
x"A8367D16",
x"A7FA7D0F",
x"A7CC7D2C",
x"A7AE7D6B",
x"A7A27DC1",
x"A7AE7E26",
x"A7CF7E8C",
x"A8087EE8",
x"A8567F2F",
x"A8B37F5D",
x"A9147F6D",
x"A96E7F60",
x"A9B57F36",
x"A9DD7EF5",
x"A9DD7E9F",
x"A9AE7E39",
x"A94F7DC4",
x"A8C27D44",
x"A80E7CBA",
x"A73C7C28",
x"A6547B8E",
x"A5627AEE",
x"A46A7A4B",
x"A37379AC",
x"A2807915",
x"A194788C",
x"A0AC7818",
x"9FCC77BA",
x"9EF07778",
x"9E1C774E",
x"9D52773A",
x"9C977736",
x"9BF1773A",
x"9B6B7741",
x"9B0E7746",
x"9AE47744",
x"9AF4773D",
x"9B407736",
x"9BC97734",
x"9C86773E",
x"9D6A775D",
x"9E637792",
x"9F5E77E1",
x"A0467846",
x"A10878BD",
x"A19A793C",
x"A1F079B7",
x"A20B7A26",
x"A1F07A78",
x"A1A17AA6",
x"A1227AA5",
x"A0747A6D",
x"9F8D79F4",
x"9E5F7934",
x"9CCF7829",
x"9AC876CE",
x"98317523",
x"94FA732D",
x"912470F5",
x"8CBE6E8D",
x"87EC6C0F",
x"82E66996",
x"7DEF6742",
x"79526537",
x"75596390",
x"72456264",
x"704461C3",
x"6F6F61B2",
x"6FC86228",
x"71386314",
x"7397645F",
x"76B065EC",
x"7A45679E",
x"7E20695C",
x"820D6B10",
x"85E96CAD",
x"899B6E2B",
x"8D1B6F89",
x"906970CE",
x"93907202",
x"969B732F",
x"999A745C",
x"9C957592",
x"9F9276D5",
x"A2927823",
x"A58D7979",
x"A8787AD0",
x"AB467C20",
x"ADE77D5E",
x"B04F7E84",
x"B2707F87",
x"B4438063",
x"B5C38115",
x"B6F3819E",
x"B7D18200",
x"B867823F",
x"B8BF8263",
x"B8E38274",
x"B8DE827A",
x"B8B9827B",
x"B87E8280",
x"B833828A",
x"B7DD829C",
x"B77B82B5",
x"B70E82D1",
x"B69682EE",
x"B6118308",
x"B57E8317",
x"B4E1831B",
x"B43C830F",
x"B39782FA",
x"B2F782DC",
x"B26A82BF",
x"B1F682A9",
x"B1A682A5",
x"B18282B9",
x"B18F82E8",
x"B1CA8335",
x"B2308395",
x"B2B68402",
x"B34C846D",
x"B3DD84C2",
x"B45484F3",
x"B49984F0",
x"B49984B2",
x"B4448436",
x"B3928382",
x"B28582A3",
x"B12881AD",
x"AF9180B6",
x"ADDE7FD7",
x"AC387F26",
x"AABF7EB5",
x"A99E7E8B",
x"A8F57EAD",
x"A8DF7F1B",
x"A9677FC9",
x"AA9280AB",
x"AC5781B0",
x"AE9E82CC",
x"B14A83ED",
x"B4338507",
x"B72F8611",
x"BA128701",
x"BCB487D4",
x"BEF48885",
x"C0BA8914",
x"C1FA8980",
x"C2AF89CA",
x"C2E489F6",
x"C2A98A04",
x"C21689FB",
x"C14489DD",
x"C04C89B1",
x"BF3D8979",
x"BE298936",
x"BD1188EE",
x"BBF488A1",
x"BACD884D",
x"B99487F6",
x"B846879D",
x"B6E48742",
x"B57B86EA",
x"B41E869B",
x"B2E78657",
x"B1F28628",
x"B160860F",
x"B143860E",
x"B1A68622",
x"B2878648",
x"B3D08678",
x"B56486A8",
x"B71B86CD",
x"B8CC86E3",
x"BA4E86E2",
x"BB8586C9",
x"BC5D869F",
x"BCD0866C",
x"BCE58638",
x"BCA6860B",
x"BC2085ED",
x"BB5885D7",
x"BA4C85C2",
x"B8ED8598",
x"B722853D",
x"B4CA8495",
x"B1C5837D",
x"ADF881DD",
x"A95B7FA6",
x"A3F77CDB",
x"9DEE798C",
x"977E75DC",
x"90F37203",
x"8AAA6E3D",
x"84FD6ACB",
x"804567E9",
x"7CC565CB",
x"7AAA648E",
x"7A00643E",
x"7AB964CC",
x"7CAD661A",
x"7F9E67FA",
x"83426A35",
x"874F6C94",
x"8B7B6EE6",
x"8F917108",
x"936272E5",
x"96D77476",
x"99EA75C7",
x"9CA176E8",
x"9F1177F4",
x"A15078FE",
x"A37D7A1D",
x"A5AC7B5D",
x"A7F87CBF",
x"AA707E3D",
x"AD1C7FCF",
x"B0028167",
x"B32182F7",
x"B66B8474",
x"B9D685D7",
x"BD49871E",
x"C0AC8848",
x"C3E18958",
x"C6CA8A4D",
x"C9478B28",
x"CB3D8BE0",
x"CC988C71",
x"CD4B8CD2",
x"CD558CF9",
x"CCC78CE3",
x"CBB78C97",
x"CA4C8C1B",
x"C8B28B88",
x"C7188AF7",
x"C5AA8A85",
x"C4918A50",
x"C3E18A6D",
x"C3A88AE9",
x"C3DA8BC3",
x"C4618CEF",
x"C51E8E4F",
x"C5E78FC4",
x"C6959127",
x"C70C9258",
x"C73D9341",
x"C72993D6",
x"C6E2941E",
x"C68E942B",
x"C657941A",
x"C66D940E",
x"C6F89428",
x"C8129480",
x"C9C39524",
x"CBFC9611",
x"CE99973A",
x"D16A9882",
x"D43699CA",
x"D6C79AF2",
x"D8F59BE4",
x"DAA69C8D",
x"DBD79CEB",
x"DC969D08",
x"DD059CF2",
x"DD4B9CC2",
x"DD939C8F",
x"DDFC9C69",
x"DE9D9C5B",
x"DF769C68",
x"E07F9C8C",
x"E1A09CBA",
x"E2BB9CE9",
x"E3B69D0F",
x"E47B9D29",
x"E4FD9D36",
x"E5409D3D",
x"E54B9D48",
x"E5319D64",
x"E5019D93",
x"E4C49DD5",
x"E4829E22",
x"E42E9E65",
x"E3BB9E86",
x"E30D9E69",
x"E2069DF5",
x"E08D9D12",
x"DE8D9BB8",
x"DBFC99EB",
x"D8DF97BA",
x"D5479542",
x"D15392AB",
x"CD26901D",
x"C8EE8DBF",
x"C4DA8BB5",
x"C1128A14",
x"BDB988E6",
x"BAE78825",
x"B8A887BC",
x"B6F78791",
x"B5C4877E",
x"B4F1875E",
x"B457870F",
x"B3C78676",
x"B3198582",
x"B2268432",
x"B0D3828A",
x"AF18809F",
x"ACFB7E8E",
x"AA927C72",
x"A7FD7A6B",
x"A5647896",
x"A2EA7703",
x"A0A675BA",
x"9EA274B7",
x"9CCC73EB",
x"9B03733B",
x"9915728A",
x"96C871B9",
x"93E370A9",
x"903E6F47",
x"8BC56D88",
x"86866B6B",
x"80AA6901",
x"7A796663",
x"745263B4",
x"6E996117",
x"69B15EB3",
x"65EE5CAB",
x"63825B15",
x"62855A01",
x"62E85975",
x"647A596A",
x"66F659D2",
x"6A065A98",
x"6D525BA6",
x"708D5CE1",
x"737A5E33",
x"75F25F87",
x"77E560CB",
x"795861F3",
x"7A5F62F6",
x"7B1863CC",
x"7BA06477",
x"7C1164F4",
x"7C7C654B",
x"7CE86580",
x"7D58659B",
x"7DC565AA",
x"7E2A65B7",
x"7E8065CB",
x"7EC865F2",
x"7F066630",
x"7F426687",
x"7F8A66F9",
x"7FE9677F",
x"80676811",
x"810D68A7",
x"81D66937",
x"82BE69BA",
x"83B56A28",
x"84B16A83",
x"859E6AC8",
x"86716AFA",
x"87216B20",
x"87A86B3B",
x"880A6B52",
x"884B6B69",
x"88746B83",
x"88906B9E",
x"88A76BBE",
x"88C36BDF",
x"88E96C00",
x"891B6C21",
x"89566C3F",
x"89976C5B",
x"89D86C72",
x"8A116C82",
x"8A3B6C8A",
x"8A4F6C87",
x"8A486C78",
x"8A226C58",
x"89E06C27",
x"89816BE2",
x"890B6B8A",
x"88836B1E",
x"87EC6A9E",
x"874D6A0F",
x"86AC696F",
x"860A68C5",
x"85666814",
x"84C16766",
x"841866C1",
x"836C6631",
x"82BC65BF",
x"820D6579",
x"81636565",
x"80CC658D",
x"805165EF",
x"8000668A",
x"7FE66753",
x"800E683B",
x"807A692E",
x"812D6A17",
x"821E6AE1",
x"83426B7C",
x"84896BDF",
x"85E06C06",
x"87356BF8",
x"88746BC1",
x"89906B72",
x"8A7C6B20",
x"8B316ADC",
x"8BAB6AB5",
x"8BE76AB1",
x"8BE96AD2",
x"8BB16B10",
x"8B426B5F",
x"8AA26BB0",
x"89D56BEF",
x"88E06C13",
x"87CC6C12",
x"86A06BE6",
x"85636B96",
x"84246B27",
x"82EC6AA8",
x"81C56A23",
x"80B869A3",
x"7FCC6931",
x"7F0468CF",
x"7E60687D",
x"7DDC6835",
x"7D6F67F0",
x"7D0D67A7",
x"7CAA6753",
x"7C3966F3",
x"7BB4668A",
x"7B11661E",
x"7A4F65BA",
x"79706568",
x"787F6535",
x"77836528",
x"76876541",
x"7597657C",
x"74B565C8",
x"73DF660E",
x"730D6634",
x"722B661B",
x"712665A8",
x"6FE264C4",
x"6E4C6360",
x"6C556181",
x"69F75F33",
x"67415C92",
x"644759C7",
x"613056FE",
x"5E29546B",
x"5B62523A",
x"590C508F",
x"574E4F86",
x"56444F25",
x"55F64F65",
x"56615033",
x"5773516D",
x"591052E8",
x"5B135481",
x"5D5B560C",
x"5FC45771",
x"6234589A",
x"64995980",
x"66E45A26",
x"690C5A9B",
x"6B0E5AF1",
x"6CE95B3C",
x"6E995B90",
x"701B5BF7",
x"716D5C7D",
x"728C5D21",
x"73735DDD",
x"74275EA7",
x"74AA5F72",
x"7502602F",
x"753760D8",
x"7552615F",
x"755C61C5",
x"75596209",
x"754C622D",
x"753A6239",
x"751D6237",
x"74F6622B",
x"74C4621E",
x"74876213",
x"7445620D",
x"74006209",
x"73C16204",
x"738E61FC",
x"736F61E9",
x"736661C6",
x"73766193",
x"739E614B",
x"73D860F3",
x"741D6091",
x"7468602B",
x"74B15FCC",
x"74F25F81",
x"752A5F50",
x"75555F42",
x"75765F5C",
x"758C5F9A",
x"759B5FF6",
x"75A56067",
x"75AE60DF",
x"75B46150",
x"75BA61AB",
x"75BC61E6",
x"75BC61FC",
x"75B761E8",
x"75A861B1",
x"758C615D",
x"755E60F7",
x"751D608D",
x"74C56029",
x"74585FD8",
x"73DB5F9D",
x"73535F7E",
x"72CC5F7D",
x"72555F9A",
x"71FC5FCD",
x"71CE6018",
x"71D66074",
x"721D60DD",
x"72A0614E",
x"735661C2",
x"74316231",
x"751B6297",
x"760062EC",
x"76C46327",
x"77536344",
x"77A1633E",
x"77A56315",
x"776062CC",
x"76DC6266",
x"762861EF",
x"7558616F",
x"747F60F0",
x"73AD607C",
x"72F36014",
x"72565FBE",
x"71DB5F76",
x"717F5F39",
x"71375F01",
x"70FC5EC8",
x"70C25E8A",
x"70815E45",
x"70355DFD",
x"6FDB5DB6",
x"6F765D78",
x"6F0F5D4B",
x"6EAA5D33",
x"6E565D35",
x"6E1A5D52",
x"6DFD5D86",
x"6E035DC9",
x"6E285E14",
x"6E665E5C",
x"6EB55E9A",
x"6F065EC5",
x"6F4C5EDA",
x"6F7A5ED7",
x"6F895EBF",
x"6F6C5E92",
x"6F245E55",
x"6EB05E0A",
x"6E105DB1",
x"6D485D4C",
x"6C5B5CD7",
x"6B4B5C50",
x"6A1A5BB6",
x"68CC5B08",
x"67645A45",
x"65E85970",
x"64625892",
x"62E157B6",
x"617656E6",
x"60355630",
x"5F3755A2",
x"5E8C5547",
x"5E43552B",
x"5E635550",
x"5EEE55BC",
x"5FD8566D",
x"6111575C",
x"62895881",
x"642859D3",
x"65E15B46",
x"67A75CD0",
x"69795E64",
x"6B595FF9",
x"6D526184",
x"6F7062FD",
x"71BE645C",
x"74416598",
x"76F266AE",
x"79C26797",
x"7C9B6852",
x"7F5D68DE",
x"81E66941",
x"841B6984",
x"85E769B5",
x"874569E3",
x"883B6A23",
x"88DF6A82",
x"89556B0F",
x"89BE6BD2",
x"8A3E6CCD",
x"8AEF6DF5",
x"8BDC6F3E",
x"8D03708F",
x"8E4F71CF",
x"8FA172E6",
x"90D873C0",
x"91D0744E",
x"9276748C",
x"92C0747F",
x"92B97436",
x"927A73C7",
x"922B734B",
x"91F672DB",
x"9205728A",
x"92777265",
x"93597274",
x"94A772B0",
x"964C7312",
x"9822738C",
x"9A01740F",
x"9BBE748F",
x"9D367505",
x"9E59756F",
x"9F2475D2",
x"9FA47636",
x"9FF176A6",
x"A031772C",
x"A08077D1",
x"A0F97896",
x"A1A67977",
x"A2887A65",
x"A3907B54",
x"A4A17C2D",
x"A59B7CDE",
x"A6607D59",
x"A6D97D94",
x"A6FD7D91",
x"A6CD7D57",
x"A6617CFB",
x"A5D77C94",
x"A5597C3C",
x"A50B7C0B",
x"A5117C16",
x"A5827C65",
x"A6667CF8",
x"A7B07DC3",
x"A9467EAF",
x"AB017F9E",
x"ACAF8077",
x"AE21811B",
x"AF2F8177",
x"AFB8817E",
x"AFAE8133",
x"AF12809F",
x"ADF77FD7",
x"AC7E7EF4",
x"AACC7E0C",
x"A90B7D39",
x"A7617C88",
x"A5EB7C01",
x"A4BB7BA0",
x"A3D07B60",
x"A3257B2D",
x"A2A47AFC",
x"A2367ABC",
x"A1C57A63",
x"A13F79ED",
x"A09B7960",
x"9FDA78C3",
x"9F0D7825",
x"9E487793",
x"9DA5771F",
x"9D3F76D1",
x"9D2976AF",
x"9D6E76B6",
x"9E0B76E1",
x"9EEC7723",
x"9FF6776C",
x"A10177B2",
x"A1E477E1",
x"A27877F5",
x"A29F77E7",
x"A24877B7",
x"A16B776B",
x"A0187709",
x"9E66769B",
x"9C737626",
x"9A6075AF",
x"984C7534",
x"964974B0",
x"94607415",
x"92877352",
x"90A97257",
x"8EAB7110",
x"8C6C6F73",
x"89CF6D7C",
x"86C56B30",
x"834C68A4",
x"7F7765F5",
x"7B6A634B",
x"775B60D2",
x"73875EB8",
x"70305D24",
x"6D8F5C32",
x"6BD35BF6",
x"6B1A5C6D",
x"6B695D8B",
x"6CB15F32",
x"6ED4613F",
x"71A46387",
x"74F065E6",
x"78846837",
x"7C316A65",
x"7FD56C5F",
x"83556E27",
x"86A56FC0",
x"89C27135",
x"8CAF7297",
x"8F7473F2",
x"921E7552",
x"94B276BC",
x"973B782C",
x"99BC799F",
x"9C387B0B",
x"9EAC7C64",
x"A1177D9F",
x"A3717EB3",
x"A5B37F95",
x"A7D38045",
x"A9C680BF",
x"AB7D8105",
x"ACED811F",
x"AE078114",
x"AEC380E8",
x"AF1F80A9",
x"AF16805E",
x"AEB3800E",
x"AE017FC2",
x"AD117F7E",
x"ABF67F45",
x"AAC67F15",
x"A9967EF0",
x"A87B7ED0",
x"A7847EB0",
x"A6B87E8F",
x"A61E7E68",
x"A5B37E3A",
x"A5747E02",
x"A5597DC3",
x"A5527D7F",
x"A5547D36",
x"A5537CEB",
x"A5427CA0",
x"A5177C56",
x"A4CD7C09",
x"A4667BBA",
x"A3E47B67",
x"A3537B0E",
x"A2C07AB3",
x"A23B7A56",
x"A1D279FE",
x"A19279B2",
x"A1857975",
x"A1AC7950",
x"A2007944",
x"A2747953",
x"A2F6797B",
x"A37179B6",
x"A3D279FB",
x"A4027A44",
x"A3FB7A89",
x"A3B97AC3",
x"A33F7AED",
x"A29E7B08",
x"A1E77B15",
x"A1357B19",
x"A09E7B1B",
x"A0367B1F",
x"A00F7B2C",
x"A0317B43",
x"A09A7B6A",
x"A1467B9F",
x"A2267BE1",
x"A32E7C30",
x"A4477C8B",
x"A5627CED",
x"A66E7D54",
x"A75D7DBC",
x"A8257E1F",
x"A8BC7E78",
x"A91F7EBD",
x"A9497EE8",
x"A93C7EF1",
x"A8F77ED4",
x"A8807E8F",
x"A7DC7E25",
x"A7127D9F",
x"A62C7D06",
x"A5337C6A",
x"A4327BDA",
x"A3327B63",
x"A23D7B0F",
x"A15D7AE4",
x"A09E7AE1",
x"A0087B04",
x"9FA87B40",
x"9F877B8E",
x"9FB17BE1",
x"A02B7C30",
x"A0F97C75",
x"A2177CAC",
x"A37B7CD6",
x"A5147CF5",
x"A6C87D0F",
x"A87A7D29",
x"AA0B7D47",
x"AB607D6D",
x"AC5C7D99",
x"ACEE7DC9",
x"AD0B7DF2",
x"ACAB7E0E",
x"ABC97E0B",
x"AA667DD6",
x"A87B7D5E",
x"A6017C8C",
x"A2EE7B50",
x"9F39799C",
x"9ADA7768",
x"95D574B7",
x"903B7196",
x"8A2F6E1D",
x"83E76A6F",
x"7DA766B4",
x"77BE631B",
x"727D5FD0",
x"6E2D5CFD",
x"6B025AC0",
x"691D592F",
x"687F584F",
x"690A581C",
x"6A8F5884",
x"6CC85970",
x"6F6F5AC0",
x"723F5C59",
x"75065E1E",
x"779D5FF9",
x"79F961DA",
x"7C1E63B8",
x"7E20658B",
x"80146752",
x"8213690A",
x"84286AB2",
x"86586C45",
x"88946DBB",
x"8AC56F0C",
x"8CCF702A",
x"8E90710A",
x"8FF271A4",
x"90E471F2",
x"916771F5",
x"918771B3",
x"9160713A",
x"9114709F",
x"90C66FF8",
x"909A6F61",
x"90AB6EEF",
x"91066EB8",
x"91AC6EC5",
x"92956F1A",
x"93A86FAE",
x"94C87070",
x"95D37148",
x"96AE721A",
x"973F72CE",
x"9777734A",
x"97527382",
x"96D5736F",
x"96117317",
x"951C7288",
x"941471D8",
x"93147120",
x"92347079",
x"918A6FF9",
x"91216FAD",
x"91016F9C",
x"91276FC4",
x"9185701C",
x"92117092",
x"92B57116",
x"935D7193",
x"93F771F9",
x"9470723D",
x"94BE7252",
x"94D6723B",
x"94B971F8",
x"94697192",
x"93F07112",
x"93597089",
x"92B67003",
x"921B6F8F",
x"91976F3A",
x"913C6F0F",
x"91176F13",
x"912C6F47",
x"917B6FAB",
x"91FD7037",
x"92A270E1",
x"9359719A",
x"94087257",
x"949E7308",
x"950473A1",
x"9532741C",
x"951E7472",
x"94CD74A1",
x"944674AD",
x"93987499",
x"92D3746A",
x"92057426",
x"913C73D1",
x"9081736E",
x"8FD672FE",
x"8F377280",
x"8E9B71F5",
x"8DF9715B",
x"8D4570B1",
x"8C736FFC",
x"8B7B6F3D",
x"8A5F6E7A",
x"891D6DBE",
x"87BE6D0F",
x"864F6C75",
x"84E06BF6",
x"83846B97",
x"824E6B59",
x"814C6B3A",
x"808E6B34",
x"801A6B41",
x"7FF36B55",
x"80136B69",
x"806F6B75",
x"80F46B70",
x"81906B59",
x"822B6B30",
x"82B16AFA",
x"83116ABF",
x"83416A89",
x"833C6A5E",
x"83046A45",
x"829E6A42",
x"82156A51",
x"81706A68",
x"80B16A79",
x"7FD66A73",
x"7ED66A41",
x"7DA369D1",
x"7C2A6914",
x"7A586804",
x"7820669E",
x"757C64ED",
x"727662FE",
x"6F2060E9",
x"6B9C5EC5",
x"68135CAC",
x"64B75AB8",
x"61BA58FA",
x"5F45577F",
x"5D7D5651",
x"5C725570",
x"5C2A54DA",
x"5C965488",
x"5D9E5473",
x"5F205494",
x"60F254E0",
x"62ED5556",
x"64EE55F0",
x"66D556A9",
x"6893577F",
x"6A1A5870",
x"6B6C5973",
x"6C8A5A81",
x"6D835B95",
x"6E5F5CA5",
x"6F2B5DA7",
x"6FF05E92",
x"70B85F63",
x"71846015",
x"725860A7",
x"732E611E",
x"7406617E",
x"74D861D3",
x"75A16222",
x"765C6276",
x"770462D3",
x"7798633E",
x"781663B7",
x"787D6437",
x"78D264B5",
x"7916652A",
x"794E6587",
x"797D65C2",
x"79A865D2",
x"79D365B2",
x"79FF6565",
x"7A2764EC",
x"7A4E6453",
x"7A6C63A8",
x"7A7D62FC",
x"7A80625F",
x"7A6F61E2",
x"7A496193",
x"7A136179",
x"79CE6198",
x"798061F0",
x"79346277",
x"78F26321",
x"78BE63DC",
x"78A16497",
x"789E653F",
x"78B865C8",
x"78EB6621",
x"79356648",
x"7990663C",
x"79F46601",
x"7A5C65A7",
x"7ABE6538",
x"7B1364C8",
x"7B536465",
x"7B77641B",
x"7B7C63F3",
x"7B5E63EC",
x"7B1B6401",
x"7AB9642B",
x"7A41645A",
x"79BB6486",
x"793464A3",
x"78BB64AA",
x"7860649E",
x"782E6484",
x"782D6469",
x"785F6459",
x"78C16463",
x"794B6493",
x"79EC64E9",
x"7A946566",
x"7B3165FF",
x"7BB166A4",
x"7C07673F",
x"7C2D67BB",
x"7C1E6806",
x"7BE06813",
x"7B7D67DE",
x"7AFE676B",
x"7A7366C5",
x"79E56604",
x"795D653E",
x"78E06489",
x"787263FA",
x"780E639F",
x"77B5637F",
x"77636395",
x"771463D9",
x"76C96439",
x"768664A4",
x"764B6504",
x"761E654C",
x"76066572",
x"7606656D",
x"761D6542",
x"764C64FA",
x"768F64A0",
x"76DC6441",
x"772B63EC",
x"777563AB",
x"77B16386",
x"77DD637D",
x"77F7638E",
x"77FF63B4",
x"77F763E2",
x"77E3640B",
x"77C46424",
x"7798641E",
x"775963EF",
x"76FD638B",
x"767762F0",
x"75B7621A",
x"74AE6107",
x"734F5FBE",
x"71935E49",
x"6F7D5CB5",
x"6D165B12",
x"6A6D5974",
x"67A057F1",
x"64CB569B",
x"62115584",
x"5F9454B8",
x"5D725440",
x"5BC4541E",
x"5A99544A",
x"59F954BD",
x"59E5556A",
x"5A4E563D",
x"5B265728",
x"5C52581C",
x"5DB8590F",
x"5F3D59F4",
x"60C55AC9",
x"623A5B85",
x"63895C2B",
x"64AA5CB8",
x"659A5D29",
x"665E5D83",
x"67005DC2",
x"678D5DE9",
x"68175DFA",
x"68A85DF8",
x"694C5DEC",
x"6A095DD9",
x"6ADC5DC8",
x"6BBF5DC3",
x"6CA75DD0",
x"6D895DF8",
x"6E595E3F",
x"6F115EA8",
x"6FAE5F32",
x"70345FD9",
x"70AA6098",
x"711A6164",
x"71936232",
x"721A62F3",
x"72B8639B",
x"736A641D",
x"742B646F",
x"74EF648A",
x"75A76472",
x"7644642A",
x"76B863C1",
x"76FC6346",
x"770E62D2",
x"76F66277",
x"76BF6248",
x"767C6250",
x"763F6294",
x"761E6310",
x"762A63B8",
x"76726479",
x"76F9653C",
x"77C465ED",
x"78C76677",
x"79F966CF",
x"7B4466F2",
x"7C9566E0",
x"7DD866A8",
x"7EF7665B",
x"7FE2660A",
x"808D65C9",
x"80F365A7",
x"811865AE",
x"810465E2",
x"80C7663C",
x"806D66B5",
x"800D6741",
x"7FB567CF",
x"7F726852",
x"7F4868BF",
x"7F38690C",
x"7F3B6932",
x"7F426930",
x"7F416904",
x"7F2468B4",
x"7EDF6845",
x"7E6967BE",
x"7DBE6725",
x"7CDF6686",
x"7BD865E6",
x"7AB46552",
x"798464D0",
x"785B646A",
x"77486424",
x"765B6403",
x"75A06406",
x"751D6428",
x"74D66466",
x"74CB64B7",
x"74F4650B",
x"754B655E",
x"75C1659E",
x"764B65C6",
x"76D965D2",
x"776065BE",
x"77D3658D",
x"782E6545",
x"786F64F0",
x"789A6495",
x"78B76444",
x"78D36404",
x"78FA63DF",
x"793763D9",
x"798D63F6",
x"79FC6431",
x"7A7A6487",
x"7AF964ED",
x"7B656559",
x"7BAB65BE",
x"7BB9660D",
x"7B86663C",
x"7B116644",
x"7A62661D",
x"798A65C8",
x"78A16546",
x"77C164A4",
x"76FD63E8",
x"7663631F",
x"75F56255",
x"75A76193",
x"756060DF",
x"75046038",
x"746F5F9D",
x"737F5F04",
x"72205E69",
x"704B5DBF",
x"6E075D00",
x"6B705C2B",
x"68B25B42",
x"66025A4D",
x"6399595F",
x"61B05887",
x"607357E0",
x"6006577F",
x"60735778",
x"61B757D9",
x"63B858A5",
x"665259D9",
x"69555B66",
x"6C8A5D32",
x"6FC25F22",
x"72CE6113",
x"758C62E4",
x"77E56479",
x"79CF65BE",
x"7B4B66A8",
x"7C65673A",
x"7D2B677C",
x"7DB26783",
x"7E10676C",
x"7E55674E",
x"7E8E6744",
x"7EC5675F",
x"7EFC67A8",
x"7F316820",
x"7F6068BB",
x"7F836968",
x"7F966A0F",
x"7F906A9A",
x"7F6F6AF5",
x"7F326B10",
x"7EDC6AE6",
x"7E706A7D",
x"7DF269DF",
x"7D696921",
x"7CDE6859",
x"7C5667A1",
x"7BDB670D",
x"7B7066B0",
x"7B1D6691",
x"7AE366B1",
x"7AC86709",
x"7ACC678A",
x"7AEF6821",
x"7B3168B8",
x"7B8E693B",
x"7C096999",
x"7C9969C7",
x"7D3E69BE",
x"7DF26986",
x"7EB06927",
x"7F7268B2",
x"8032683C",
x"80E967D8",
x"818E6797",
x"821D6787",
x"828E67AE",
x"82DC680C",
x"83066896",
x"830B693E",
x"82EF69F0",
x"82B46A9C",
x"82636B2B",
x"82016B92",
x"81986BC7",
x"81316BCA",
x"80D16BA1",
x"807E6B5B",
x"80416B03",
x"801D6AAD",
x"80146A65",
x"802A6A3A",
x"805F6A2D",
x"80AF6A3F",
x"811B6A68",
x"81986A9C",
x"82246AC9",
x"82B16AE5",
x"83386AE1",
x"83AF6AB4",
x"84116A5E",
x"845969E2",
x"8486694B",
x"849568A7",
x"848E6806",
x"8474677A",
x"844E6711",
x"842066D5",
x"83EF66CB",
x"83BC66F2",
x"83906744",
x"836A67B8",
x"834F6841",
x"834268D4",
x"83496965",
x"836969EC",
x"83A46A63",
x"83FA6AC9",
x"84696B1D",
x"84EA6B61",
x"85736B96",
x"85F66BBF",
x"86656BE2",
x"86B56BFC",
x"86DF6C10",
x"86E06C1E",
x"86B96C24",
x"86776C24",
x"86276C1D",
x"85D56C0D",
x"85936BF5",
x"856A6BD5",
x"85636BB1",
x"857B6B89",
x"85AE6B61",
x"85EF6B3B",
x"862E6B1D",
x"86596B07",
x"865D6AF9",
x"86276AED",
x"85A16ADC",
x"84BA6AB5",
x"835D6A68",
x"817E69DC",
x"7F0E68FF",
x"7C0A67BB",
x"78726607",
x"745663E2",
x"6FD46156",
x"6B135E7E",
x"664E5B80",
x"61C15885",
x"5DB055C3",
x"5A585366",
x"57EE5198",
x"568F5071",
x"56434FFC",
x"56FB5033",
x"588C50FC",
x"5ABE5237",
x"5D4B53B9",
x"5FE95556",
x"625B56E7",
x"646D5850",
x"66035981",
x"67145A74",
x"67AD5B32",
x"67EB5BC9",
x"67F25C4C",
x"67EE5CCB",
x"68005D52",
x"68425DE6",
x"68C15E86",
x"697C5F25",
x"6A665FB9",
x"6B6C602F",
x"6C75607A",
x"6D6C6093",
x"6E3F6076",
x"6EE56029",
x"6F5B5FB8",
x"6FA35F35",
x"6FC65EB1",
x"6FD45E41",
x"6FD45DF3",
x"6FD25DD5",
x"6FD45DE9",
x"6FDE5E2E",
x"6FED5E9E",
x"70055F2E",
x"701D5FD0",
x"70356074",
x"704E610B",
x"7068618D",
x"708961EF",
x"70B5622E",
x"70F6624F",
x"71586258",
x"71E26258",
x"729D6259",
x"738E626D",
x"74BA62A2",
x"761A62FE",
x"77A76386",
x"79526432",
x"7B0964F9",
x"7CB565C6",
x"7E3F6689",
x"7F936728",
x"809E6794",
x"815567C4",
x"81B967B4",
x"81D06770",
x"81AE6709",
x"816A6696",
x"81226634",
x"80F365FD",
x"80F66604",
x"813E6656",
x"81D366F5",
x"82B567D3",
x"83D568E3",
x"851D6A0C",
x"86736B31",
x"87B76C41",
x"88CF6D26",
x"89A56DD8",
x"8A2B6E55",
x"8A5D6EA1",
x"8A426EC5",
x"89E36ECF",
x"89566ECA",
x"88AB6EBF",
x"87F66EB5",
x"87466EAD",
x"86A56EA6",
x"86176E9C",
x"859A6E88",
x"85276E65",
x"84BB6E31",
x"84506DEE",
x"83E36D9A",
x"83736D3B",
x"83036CD4",
x"82986C69",
x"82356BFD",
x"81DF6B90",
x"81936B20",
x"814B6AAA",
x"81006A2A",
x"80A4699A",
x"802B68F9",
x"7F896845",
x"7EB5677F",
x"7DAF66AB",
x"7C7A65D0",
x"7B2564F6",
x"79BE6424",
x"78596365",
x"770B62BF",
x"75E8623B",
x"74FA61DA",
x"744C61A1",
x"73DC618E",
x"73A3619D",
x"739361C9",
x"739D6207",
x"73AD624F",
x"73AB6291",
x"738462C2",
x"732462CF",
x"727A62AD",
x"717A624F",
x"701A61A9",
x"6E5860BC",
x"6C375F86",
x"69C55E0E",
x"67145C64",
x"64445A9B",
x"617258CC",
x"5ECA570C",
x"5C71557A",
x"5A8C5429",
x"593D532C",
x"5893528F",
x"589C5256",
x"594E527F",
x"5A975304",
x"5C5B53D3",
x"5E7654DE",
x"60C25612",
x"631A575D",
x"656158AE",
x"677F59F8",
x"696D5B33",
x"6B2A5C57",
x"6CBE5D64",
x"6E375E5D",
x"6FA55F45",
x"71196021",
x"729760F9",
x"742461CE",
x"75BB62A4",
x"7752637C",
x"78DC6453",
x"7A496525",
x"7B9065EC",
x"7CA566A3",
x"7D8A6744",
x"7E4267CB",
x"7EDC6838",
x"7F65688D",
x"7FEF68CF",
x"80876906",
x"813C693B",
x"82146979",
x"831069C7",
x"842B6A2A",
x"855D6AA6",
x"869B6B37",
x"87D96BD7",
x"890B6C7D",
x"8A2C6D1E",
x"8B356DB0",
x"8C256E26",
x"8CFB6E7A",
x"8DBB6EAA",
x"8E656EB5",
x"8EF96EA3",
x"8F7A6E7A",
x"8FE46E45",
x"903B6E12",
x"90796DE9",
x"90A26DD5",
x"90B66DD9",
x"90BB6DFA",
x"90B46E33",
x"90A86E7D",
x"909E6ED1",
x"909A6F26",
x"909F6F6C",
x"90AF6F9F",
x"90CB6FB1",
x"90EE6FA1",
x"91186F6B",
x"91466F10",
x"91766E96",
x"91A46E09",
x"91D06D72",
x"91FA6CE2",
x"921E6C68",
x"92396C10",
x"92456BE6",
x"92396BF0",
x"92136C30",
x"91C96C9E",
x"915A6D34",
x"90CB6DE1",
x"901F6E94",
x"8F666F3D",
x"8EAC6FCD",
x"8E067039",
x"8D807078",
x"8D277089",
x"8CFE7070",
x"8D047035",
x"8D2E6FDE",
x"8D6A6F73",
x"8DA56EFA",
x"8DCB6E7A",
x"8DCC6DF0",
x"8D9C6D61",
x"8D3E6CC8",
x"8CB66C28",
x"8C156B87",
x"8B716AED",
x"8ADF6A65",
x"8A7369FD",
x"8A3F69C7",
x"8A5069CE",
x"8AA56A19",
x"8B3B6AAA",
x"8C036B7A",
x"8CF06C7A",
x"8DE96D94",
x"8EDA6EAE",
x"8FAC6FAE",
x"904D707E",
x"90AE7108",
x"90C37145",
x"908A7134",
x"900670DF",
x"8F417052",
x"8E496FA4",
x"8D356EE8",
x"8C1A6E30",
x"8B0D6D8A",
x"8A1A6CFD",
x"894B6C84",
x"88976C17",
x"87ED6BA6",
x"872F6B19",
x"86366A5B",
x"84D66954",
x"82E867F7",
x"8048663A",
x"7CE86420",
x"78C961B2",
x"74065F08",
x"6ECC5C42",
x"695C5981",
x"640356EE",
x"5F1054AC",
x"5ACE52DA",
x"577C518F",
x"554050D7",
x"542E50AD",
x"54405107",
x"555451CD",
x"573B52E1",
x"59B85423",
x"5C8C5577",
x"5F7856BF",
x"624557E7",
x"64CF58E7",
x"66FF59BC",
x"68CE5A6B",
x"6A415B01",
x"6B695B8B",
x"6C5C5C18",
x"6D305CB3",
x"6DF85D66",
x"6EC15E2E",
x"6F935F07",
x"706D5FE4",
x"714960B9",
x"721E6174",
x"72E26206",
x"73896263",
x"740E6286",
x"746F6270",
x"74AD6228",
x"74CF61BF",
x"74DC6145",
x"74DF60CE",
x"74E3606D",
x"74EF6031",
x"75096022",
x"75326042",
x"756A608D",
x"75AE60F9",
x"75F66176",
x"763B61F6",
x"7676626F",
x"76A462D5",
x"76C16323",
x"76CE635C",
x"76D16383",
x"76CC639F",
x"76CB63B8",
x"76D463D3",
x"76EF63F6",
x"7721641D",
x"776F6448",
x"77DB6473",
x"78626498",
x"78FF64B4",
x"79AE64C4",
x"7A6664C9",
x"7B1E64C6",
x"7BCC64C1",
x"7C6664BE",
x"7CDF64BF",
x"7D3164CB",
x"7D5364DF",
x"7D4464FC",
x"7D03651E",
x"7C996542",
x"7C146565",
x"7B876587",
x"7B0965A8",
x"7AB265CE",
x"7A9B65FC",
x"7AD26638",
x"7B636684",
x"7C4B66E6",
x"7D7A6759",
x"7EDB67DB",
x"80496860",
x"81A468DE",
x"82C56948",
x"838E6990",
x"83ED69AD",
x"83DA6997",
x"835D6948",
x"828A68C5",
x"81796811",
x"804E673B",
x"7F24664E",
x"7E18655E",
x"7D3C647C",
x"7C9963B9",
x"7C2E6325",
x"7BF362C9",
x"7BDB62AA",
x"7BD862C6",
x"7BDB6318",
x"7BDC6393",
x"7BD36425",
x"7BC164BF",
x"7BA46550",
x"7B8465C8",
x"7B63661E",
x"7B45664C",
x"7B2A6653",
x"7B10663A",
x"7AF76604",
x"7ADC65C2",
x"7ABB657A",
x"7A916537",
x"7A5F64FF",
x"7A2564D5",
x"79E964B7",
x"79AD64A4",
x"79756495",
x"79486487",
x"792A6476",
x"791A645C",
x"791B643B",
x"7925640E",
x"793463D8",
x"79376393",
x"791E633E",
x"78D562D2",
x"78446249",
x"7756619E",
x"75F960CC",
x"74215FCC",
x"71CC5EA4",
x"6F045D57",
x"6BE25BF1",
x"68895A84",
x"65265922",
x"61EB57DF",
x"5F0D56D0",
x"5CBA5605",
x"5B135589",
x"5A305563",
x"5A105591",
x"5AA95608",
x"5BDE56BF",
x"5D8557A4",
x"5F7258A5",
x"617B59AF",
x"63725AB6",
x"653E5BAC",
x"66CB5C87",
x"68145D45",
x"69215DE2",
x"69FF5E60",
x"6AC45EC3",
x"6B845F10",
x"6C565F4D",
x"6D485F80",
x"6E5F5FAE",
x"6F9A5FDC",
x"70F3600E",
x"725B6049",
x"73C1608E",
x"751160DD",
x"763F6137",
x"773E6197",
x"780761FE",
x"789B6268",
x"790362D2",
x"79486339",
x"797A639D",
x"79A863FC",
x"79E26456",
x"7A3164AE",
x"7A9D6500",
x"7B286550",
x"7BD1659E",
x"7C9065E6",
x"7D5F6625",
x"7E35665B",
x"7F0B6680",
x"7FD86694",
x"80976694",
x"81456683",
x"81E06666",
x"82666646",
x"82D96630",
x"833E6632",
x"8394665F",
x"83E566C1",
x"84346763",
x"84846849",
x"84DC696C",
x"853E6ABD",
x"85A56C26",
x"860E6D88",
x"86706EC4",
x"86C16FBD",
x"86F77058",
x"87077089",
x"86EF704D",
x"86AE6FB0",
x"864C6ECB",
x"85D96DBF",
x"85696CB4",
x"85116BCC",
x"84E66B2A",
x"84FA6AE1",
x"85566AF6",
x"85F96B66",
x"86D96C1A",
x"87E66CF9",
x"89066DE2",
x"8A1E6EB8",
x"8B146F64",
x"8BD36FD4",
x"8C4B7006",
x"8C777002",
x"8C596FD5",
x"8BFD6F92",
x"8B736F4A",
x"8AD06F0D",
x"8A2B6EE4",
x"89986ECF",
x"89286ECB",
x"88E46EC7",
x"88D06EB7",
x"88E66E8D",
x"89186E3F",
x"89566DCA",
x"898A6D31",
x"899E6C83",
x"89816BD4",
x"892D6B3B",
x"88A16ACF",
x"87EC6AAA",
x"87256AD9",
x"86716B65",
x"85F46C4E",
x"85D26D88",
x"862A6EFE",
x"870B7097",
x"88777237",
x"8A5D73BE",
x"8C9B7510",
x"8F067617",
x"916A76C6",
x"93977713",
x"95627705",
x"96AB76A2",
x"976475FB",
x"978B7521",
x"9729742C",
x"96507326",
x"9511721F",
x"937D711C",
x"919E701D",
x"8F776F1E",
x"8D066E17",
x"8A456CFC",
x"872C6BC4",
x"83C16A69",
x"800968EB",
x"7C1A674B",
x"78146597",
x"742063DA",
x"706B6227",
x"6D20608E",
x"6A655F21",
x"68585DE9",
x"67045CED",
x"66685C31",
x"66735BB1",
x"67095B64",
x"68055B47",
x"69415B50",
x"6A9A5B78",
x"6BF35BBB",
x"6D385C17",
x"6E5E5C8A",
x"6F685D12",
x"705B5DAF",
x"71455E5C",
x"72355F14",
x"73325FCF",
x"74456086",
x"7569612F",
x"769961C3",
x"77C56241",
x"78E062A7",
x"79DD62F9",
x"7AB2633F",
x"7B5F6384",
x"7BE963D5",
x"7C5E6439",
x"7CCE64BB",
x"7D4C655C",
x"7DE8661A",
x"7EA766EC",
x"7F8667C6",
x"80746899",
x"815C694F",
x"821869D9",
x"82876A24",
x"82896A27",
x"820969DC",
x"81006945",
x"7F766869",
x"7D896759",
x"7B5E662B",
x"792864F4",
x"771B63CE",
x"756962D0",
x"7435620E",
x"73976195",
x"73966170",
x"7425619E",
x"752D621B",
x"768962DF",
x"781463D8",
x"79A864F7",
x"7B27662D",
x"7C776765",
x"7D906891",
x"7E6C69A6",
x"7F0E6A93",
x"7F806B55",
x"7FC86BE2",
x"7FF06C3B",
x"7FFC6C5F",
x"7FF06C51",
x"7FCF6C19",
x"7F9B6BBE",
x"7F5B6B4F",
x"7F186AD8",
x"7EE06A69",
x"7EC46A0D",
x"7ED269D1",
x"7F1769BA",
x"7F9A69CB",
x"80596A02",
x"81496A58",
x"82596AC4",
x"83706B38",
x"84746BAB",
x"85526C12",
x"85FD6C65",
x"86736CA4",
x"86BC6CCD",
x"86F06CE5",
x"87276CF0",
x"877C6CF8",
x"88076CFF",
x"88D56D0A",
x"89E26D1A",
x"8B226D2E",
x"8C766D44",
x"8DBB6D58",
x"8EC56D63",
x"8F746D65",
x"8FA96D59",
x"8F5C6D3F",
x"8E8D6D16",
x"8D506CDE",
x"8BC86C99",
x"8A1A6C48",
x"88726BED",
x"86F76B89",
x"85C96B1C",
x"84FB6AA7",
x"84916A2E",
x"848369B1",
x"84BB6937",
x"852068C1",
x"85916856",
x"85F367F9",
x"862E67AD",
x"86316775",
x"85F76751",
x"85896745",
x"84F3674E",
x"844C676B",
x"83AB679B",
x"832767D9",
x"82CE6820",
x"82A16868",
x"829868A3",
x"829E68C7",
x"829168C4",
x"8249688A",
x"819D680D",
x"80696742",
x"7E966625",
x"7C1D64BB",
x"790C630D",
x"7583612E",
x"71B15F37",
x"6DD55D45",
x"6A305B76",
x"66FD59EA",
x"647558B8",
x"62BA57F1",
x"61E1579F",
x"61E957C5",
x"62C25854",
x"644B5940",
x"665E5A6E",
x"68CB5BC8",
x"6B695D2F",
x"6E115E8E",
x"70A45FCF",
x"730E60E6",
x"754461CF",
x"7741628B",
x"790A6328",
x"7AA863AF",
x"7C256437",
x"7D8E64CC",
x"7EEC657F",
x"80486656",
x"81A56751",
x"8304686B",
x"84636997",
x"85BC6AC2",
x"87076BDC",
x"883E6CD2",
x"89566D97",
x"8A4F6E23",
x"8B246E76",
x"8BD56E94",
x"8C696E8A",
x"8CE56E66",
x"8D536E3A",
x"8DBE6E0F",
x"8E2C6DF3",
x"8EA56DEC",
x"8F296DF9",
x"8FB96E1A",
x"904F6E4A",
x"90E46E86",
x"91736EC8",
x"91F46F13",
x"92646F66",
x"92C86FCA",
x"93257040",
x"938B70D2",
x"940D7186",
x"94BE725C",
x"95AF7354",
x"96F17464",
x"988A7583",
x"9A7476A0",
x"9C9C77A9",
x"9EE6788C",
x"A126793A",
x"A33279A3",
x"A4D979C3",
x"A5F07998",
x"A65A7928",
x"A60B7881",
x"A50B77B4",
x"A37676D8",
x"A1777603",
x"9F4C754A",
x"9D3274BB",
x"9B667462",
x"9A177441",
x"99607452",
x"994A7489",
x"99C274D7",
x"9A9F752A",
x"9BB1756E",
x"9CBC7597",
x"9D88759D",
x"9DED757F",
x"9DD37543",
x"9D3974F4",
x"9C3574A0",
x"9AEF7458",
x"9997742C",
x"98627421",
x"977A743D",
x"97007478",
x"96FD74C7",
x"97647516",
x"98187550",
x"98E97561",
x"99A27534",
x"9A0E74BE",
x"9A0173FC",
x"996072F4",
x"982271B3",
x"96557051",
x"94176EEC",
x"91956DA3",
x"8F046C94",
x"8C9B6BD8",
x"8A8B6B7D",
x"88F96B8D",
x"87FA6BFF",
x"87966CC4",
x"87C26DC2",
x"88666EDE",
x"89606FF0",
x"8A8B70DE",
x"8BBC718C",
x"8CCD71E8",
x"8DA471EB",
x"8E2A7199",
x"8E5570FC",
x"8E257029",
x"8DA46F34",
x"8CE06E33",
x"8BEA6D3A",
x"8AD56C55",
x"89A96B89",
x"886D6AD4",
x"871D6A2B",
x"85AA6982",
x"840668C4",
x"821A67E3",
x"7FD366D2",
x"7D28658B",
x"7A17640E",
x"76AD6263",
x"7304609D",
x"6F475ED0",
x"6BA35D1A",
x"684E5B91",
x"65795A50",
x"634E5969",
x"61E558E7",
x"614758CD",
x"616B5914",
x"623659AC",
x"63855A82",
x"652A5B80",
x"66FC5C8A",
x"68D25D8B",
x"6A905E74",
x"6C245F3B",
x"6D8A5FDC",
x"6EC46059",
x"6FDC60BC",
x"70E1610E",
x"71DC6159",
x"72D661A7",
x"73D261FC",
x"74CB6256",
x"75BA62B7",
x"76966314",
x"77526368",
x"77EC63AA",
x"785D63D6",
x"78AA63EC",
x"78D863EC",
x"78F363DA",
x"790963BF",
x"792463A5",
x"79526391",
x"7998638D",
x"79FC639A",
x"7A7D63BB",
x"7B1763EF",
x"7BC26434",
x"7C776484",
x"7D2A64DF",
x"7DD06541",
x"7E6365A5",
x"7EDD660E",
x"7F3C667A",
x"7F8066E8",
x"7FAC6755",
x"7FCB67C2",
x"7FE2682A",
x"7FFC688A",
x"802568DE",
x"80666921",
x"80C26954",
x"813C6975",
x"81D3698A",
x"82816996",
x"834269A3",
x"840B69B5",
x"84D569D8",
x"859A6A0F",
x"86566A5C",
x"87086AC2",
x"87B46B3B",
x"885A6BC2",
x"89036C4F",
x"89B16CD9",
x"8A636D59",
x"8B1A6DCD",
x"8BCF6E2D",
x"8C7A6E7D",
x"8D106EC1",
x"8D876EFE",
x"8DD56F38",
x"8DF36F75",
x"8DDF6FB7",
x"8D986FFF",
x"8D277047",
x"8C937086",
x"8BE670B4",
x"8B2C70C3",
x"8A7070A9",
x"89B9705A",
x"89086FD2",
x"88606F13",
x"87BF6E21",
x"87206D0A",
x"86806BE1",
x"85DD6AB5",
x"853B699E",
x"849D68B0",
x"840767F7",
x"8386677D",
x"831E6746",
x"82DA674F",
x"82BC678E",
x"82C267F9",
x"82E96881",
x"8327691A",
x"837269BB",
x"83BF6A5E",
x"840A6B00",
x"844E6BA1",
x"848B6C44",
x"84CB6CE9",
x"85156D90",
x"85746E34",
x"85F06ECE",
x"868B6F58",
x"87456FC5",
x"8813700F",
x"88E47031",
x"89A5702B",
x"8A417003",
x"8AA56FC4",
x"8AC26F7A",
x"8A906F33",
x"8A0D6EF6",
x"893C6ECA",
x"88246EA7",
x"86CC6E85",
x"853C6E4E",
x"837A6DEC",
x"81876D48",
x"7F666C54",
x"7D1A6B03",
x"7AA8695B",
x"7821676D",
x"75996555",
x"732A6339",
x"70FA6146",
x"6F2D5FA5",
x"6DE55E7D",
x"6D3F5DE6",
x"6D545DF0",
x"6E285E9D",
x"6FBC5FDD",
x"7204619B",
x"74EA63B9",
x"78586617",
x"7C2E6891",
x"80536B0F",
x"84AE6D76",
x"89276FB9",
x"8DA871CD",
x"922273B0",
x"96817565",
x"9ABB76F1",
x"9EC0785D",
x"A28B79B2",
x"A6177AF7",
x"A9617C32",
x"AC707D6A",
x"AF467EA0",
x"B1EE7FD0",
x"B46A80FA",
x"B6BA8214",
x"B8DA8317",
x"BABF83FA",
x"BC5E84B8",
x"BDAA854C",
x"BE9C85BB",
x"BF30860A",
x"BF728646",
x"BF758680",
x"BF5A86C9",
x"BF468733",
x"BF6387CA",
x"BFD48895",
x"C0B58991",
x"C20C8AB2",
x"C3D98BE3",
x"C5FF8D0B",
x"C85A8E0E",
x"CABA8ED5",
x"CCEE8F49",
x"CECA8F65",
x"D02D8F27",
x"D1058E9D",
x"D1518DDD",
x"D1228D07",
x"D0928C36",
x"CFC78B87",
x"CEE78B10",
x"CE108AD9",
x"CD5A8AE6",
x"CCCE8B2B",
x"CC6A8B93",
x"CC1F8C08",
x"CBD88C73",
x"CB7B8CBC",
x"CAF18CD5",
x"CA288CB5",
x"C9188C5D",
x"C7C18BD8",
x"C6328B32",
x"C4828A80",
x"C2CD89D6",
x"C1358946",
x"BFD788E0",
x"BED088B1",
x"BE3388BE",
x"BE098908",
x"BE54898B",
x"BF068A3C",
x"C00F8B0D",
x"C1548BEC",
x"C2B68CC5",
x"C4158D87",
x"C5508E1E",
x"C64B8E7E",
x"C6F28E9B",
x"C7338E73",
x"C7048E07",
x"C6658D5F",
x"C55D8C86",
x"C3F28B85",
x"C2368A6C",
x"C0338940",
x"BDFA8807",
x"BB9586C2",
x"B911856E",
x"B6738407",
x"B3C2828A",
x"B10480F5",
x"AE3F7F4F",
x"AB7D7D9E",
x"A8C57BF2",
x"A6287A60",
x"A3B678FB",
x"A18077D8",
x"9F977705",
x"9E08768C",
x"9CDC766B",
x"9C127699",
x"9BA57702",
x"9B85778F",
x"9B9E7826",
x"9BD578A9",
x"9C0E7901",
x"9C2E7919",
x"9C1A78EA",
x"9BBF786D",
x"9B1477A9",
x"9A1476AA",
x"98C37582",
x"972B7443",
x"955C72FE",
x"936371C3",
x"9150709A",
x"8F2C6F86",
x"8CFA6E80",
x"8AB56D7F",
x"88526C70",
x"85C26B3F",
x"82F469D9",
x"7FD5682E",
x"7C5C6634",
x"788463EC",
x"7459615F",
x"6FED5EA1",
x"6B625BD0",
x"66E2590C",
x"62A0567E",
x"5ECA5449",
x"5B905289",
x"59175157",
x"577850BC",
x"56BD50B6",
x"56DE513C",
x"57C75235",
x"59555388",
x"5B615515",
x"5DBA56BC",
x"60335863",
x"62A059F3",
x"64DF5B5A",
x"66D55C90",
x"68735D92",
x"69B45E63",
x"6A9C5F08",
x"6B355F8D",
x"6B925FF7",
x"6BC26052",
x"6BD960A2",
x"6BEC60ED",
x"6C066137",
x"6C35617D",
x"6C8061BF",
x"6CEC61F7",
x"6D7A6225",
x"6E286242",
x"6EF2624E",
x"6FCE6245",
x"70B7622B",
x"719E6203",
x"727761D3",
x"733A61A1",
x"73D66176",
x"74446159",
x"747C614F",
x"747F6159",
x"744E617A",
x"73F461AB",
x"737F61E9",
x"7300622D",
x"728C6272",
x"723462B1",
x"720762EC",
x"720E6321",
x"724C6350",
x"72BB637F",
x"734C63AB",
x"73F263D9",
x"74946404",
x"7524642A",
x"758D6444",
x"75C8644B",
x"75D16439",
x"75AB640B",
x"756563C4",
x"750D6363",
x"74B562F4",
x"74726284",
x"744F621B",
x"745961C8",
x"74946191",
x"74FA617E",
x"7583618E",
x"761E61BC",
x"76BB6201",
x"77456252",
x"77AB62A2",
x"77DF62E8",
x"77DB631A",
x"779B6332",
x"7727632D",
x"7689630B",
x"75D262CF",
x"7516627C",
x"74696217",
x"73DF61AB",
x"7384613C",
x"736360D5",
x"737D607C",
x"73CE6038",
x"7449600E",
x"74E26006",
x"7583601B",
x"761B604D",
x"769B6097",
x"76F560F0",
x"7724614E",
x"772361A5",
x"76F661EC",
x"76A46218",
x"76346228",
x"75AE6218",
x"751D61ED",
x"748761AD",
x"73F6615C",
x"73706107",
x"72FA60B4",
x"729B6067",
x"72586022",
x"72325FE4",
x"72305FAC",
x"724C5F76",
x"72835F3B",
x"72CC5EFD",
x"731B5EBC",
x"73605E7C",
x"738D5E43",
x"73945E1C",
x"736C5E11",
x"73135E28",
x"72875E63",
x"71D65EC3",
x"71095F3F",
x"70315FCB",
x"6F5B6052",
x"6E9060C3",
x"6DD96108",
x"6D336114",
x"6C9660D8",
x"6BF6604F",
x"6B445F80",
x"6A735E76",
x"69765D3F",
x"68485BF4",
x"66EC5AA9",
x"656B5975",
x"63D1586A",
x"62365791",
x"60B056F3",
x"5F54568F",
x"5E3A5664",
x"5D70566A",
x"5D085698",
x"5D0556EA",
x"5D6B575A",
x"5E3757E1",
x"5F645881",
x"60E85936",
x"62B85A00",
x"64C85ADF",
x"670A5BCD",
x"69735CC8",
x"6BF55DC8",
x"6E835EC5",
x"71175FB9",
x"73A5609F",
x"76286174",
x"789A6239",
x"7AF662F2",
x"7D3563A4",
x"7F566459",
x"81516518",
x"832365E8",
x"84C466C9",
x"862F67BC",
x"876568B8",
x"885F69B2",
x"891E6AA0",
x"89A76B70",
x"89FC6C1A",
x"8A246C93",
x"8A256CD8",
x"8A046CE9",
x"89C86CCE",
x"89736C8F",
x"89086C38",
x"88886BD7",
x"87F46B73",
x"874F6B17",
x"869A6AC9",
x"85D96A8C",
x"85146A5C",
x"84556A3B",
x"83A26A24",
x"83066A14",
x"828A6A0A",
x"82326A03",
x"820669FD",
x"820469F9",
x"822D69F3",
x"827E69EC",
x"82F369E1",
x"838469CF",
x"842C69B7",
x"84E26997",
x"859B6970",
x"864E6944",
x"86EF6913",
x"877668E5",
x"87DC68BC",
x"881D689D",
x"8835688C",
x"882E688D",
x"881168A0",
x"87ED68C8",
x"87D26903",
x"87D56952",
x"880069B1",
x"88606A1E",
x"88F36A97",
x"89B46B14",
x"8A936B93",
x"8B7B6C0F",
x"8C596C82",
x"8D126CE9",
x"8D9C6D44",
x"8DED6D8D",
x"8E076DCA",
x"8DF46DF8",
x"8DC66E1C",
x"8D946E38",
x"8D706E51",
x"8D6D6E68",
x"8D956E7D",
x"8DE76E94",
x"8E5C6EAB",
x"8EE36EC1",
x"8F676ED4",
x"8FD36EE5",
x"90146EF0",
x"901E6EF8",
x"8FEE6EF8",
x"8F886EF0",
x"8EFA6EDF",
x"8E566EC5",
x"8DB56EA0",
x"8D2C6E72",
x"8CD26E3F",
x"8CB46E10",
x"8CDC6DEB",
x"8D4C6DDB",
x"8DFC6DEC",
x"8EE06E27",
x"8FE46E92",
x"90F36F29",
x"91F16FE4",
x"92C870B1",
x"9362717E",
x"93AC722B",
x"939E72A4",
x"933472D1",
x"927172A3",
x"91647217",
x"901B7134",
x"8EA87008",
x"8D1B6EA6",
x"8B7B6D26",
x"89CC6B99",
x"88036A0D",
x"86096881",
x"83C566F3",
x"81176552",
x"7DE6638D",
x"7A216193",
x"75C45F5C",
x"70E15CE6",
x"6B9C5A42",
x"662B578A",
x"60D654E4",
x"5BE5527A",
x"57A15074",
x"54474EF8",
x"51FE4E1B",
x"50DB4DE2",
x"50D84E44",
x"51D74F27",
x"53A7506A",
x"561351E1",
x"58DB5367",
x"5BC854DC",
x"5EAA5629",
x"61625745",
x"63DB5833",
x"660D58FD",
x"67FC59B3",
x"69AD5A64",
x"6B2B5B1E",
x"6C805BE6",
x"6DAF5CBD",
x"6EBE5D9F",
x"6FAD5E80",
x"707C5F53",
x"712B600E",
x"71BF60AD",
x"723A612B",
x"72A1618D",
x"72FC61DC",
x"734C621E",
x"7398625D",
x"73E062A1",
x"742462E8",
x"74636331",
x"749D6374",
x"74D263AA",
x"750363C9",
x"753763CE",
x"757063B5",
x"75B76381",
x"760B633B",
x"767262ED",
x"76E662A8",
x"77636274",
x"77E3625D",
x"785B626A",
x"78C26298",
x"791662E3",
x"79536346",
x"798063B7",
x"79A2642D",
x"79C864A1",
x"79FA6511",
x"7A44657C",
x"7AAB65E5",
x"7B316650",
x"7BD166C4",
x"7C816741",
x"7D3567C6",
x"7DDF6852",
x"7E7368DC",
x"7EE9695E",
x"7F3C69CE",
x"7F736A24",
x"7F946A5E",
x"7FAC6A79",
x"7FCB6A7A",
x"7FFC6A69",
x"804E6A51",
x"80C76A3D",
x"81686A38",
x"822F6A4C",
x"83156A80",
x"84106AD4",
x"85136B47",
x"86106BD1",
x"86FE6C6B",
x"87D56D08",
x"88906D9C",
x"89296E1C",
x"89A56E7D",
x"8A016EB8",
x"8A426EC8",
x"8A6A6EA9",
x"8A7C6E5E",
x"8A796DEE",
x"8A626D5F",
x"8A386CC1",
x"89FC6C20",
x"89AB6B89",
x"89466B0A",
x"88CF6AAD",
x"88466A77",
x"87AE6A69",
x"87086A7D",
x"865F6AAB",
x"85B56AE9",
x"85186B2B",
x"84916B69",
x"842C6B9D",
x"83F66BC7",
x"83F46BE6",
x"842F6C03",
x"84A76C24",
x"85556C4F",
x"862B6C89",
x"871B6CD1",
x"880D6D23",
x"88EC6D76",
x"89A16DC2",
x"8A1F6DFD",
x"8A5F6E1E",
x"8A5D6E24",
x"8A246E0F",
x"89BF6DE1",
x"893C6DA0",
x"88A86D52",
x"880A6CFA",
x"875F6C94",
x"869B6C19",
x"85AB6B79",
x"84746AA4",
x"82E0698C",
x"80D96826",
x"7E5B666D",
x"7B6C646D",
x"782A6238",
x"74BF5FED",
x"71665DB2",
x"6E5C5BB3",
x"6BDF5A18",
x"6A2358FE",
x"6947587D",
x"69565897",
x"6A485945",
x"6BF85A70",
x"6E355BF6",
x"70C45DB2",
x"736A5F7E",
x"75F56137",
x"783B62C1",
x"7A2D640B",
x"7BC56513",
x"7D1965DB",
x"7E3F666F",
x"7F5B66E5",
x"808E6751",
x"81F367C8",
x"8398685E",
x"85806921",
x"87A26A17",
x"89ED6B44",
x"8C456CA1",
x"8E906E24",
x"90B46FC0",
x"929E715F",
x"944572F4",
x"95A4746A",
x"96BF75B3",
x"97A576C4",
x"9860779B",
x"99017834",
x"99977896",
x"9A2B78CD",
x"9AC678E1",
x"9B6D78E2",
x"9C1E78DD",
x"9CDC78DA",
x"9DA278E2",
x"9E7078F9",
x"9F3F791F",
x"A00F7950",
x"A0DD7988",
x"A1A579C3",
x"A26479FC",
x"A31B7A36",
x"A3C97A71",
x"A46E7AAF",
x"A50F7AF7",
x"A5B27B4D",
x"A6607BB9",
x"A7227C39",
x"A8017CD0",
x"A9047D77",
x"AA2F7E25",
x"AB817ED3",
x"ACEE7F75",
x"AE698002",
x"AFDF8077",
x"B13680CD",
x"B256810A",
x"B3288130",
x"B39C814C",
x"B3A98161",
x"B350817B",
x"B29C819C",
x"B1A381C5",
x"B08181F1",
x"AF59821C",
x"AE49823D",
x"AD70824D",
x"ACE6824A",
x"ACB28232",
x"ACD68208",
x"AD4381D4",
x"ADE6819F",
x"AE9F8172",
x"AF4C8154",
x"AFCF8147",
x"B00B8147",
x"AFF38150",
x"AF7F8156",
x"AEB9814C",
x"ADAF812B",
x"AC7B80EB",
x"AB3B808F",
x"AA048019",
x"A8F07F96",
x"A8047F0F",
x"A7427E94",
x"A69F7E26",
x"A6057DCD",
x"A55E7D82",
x"A4917D3A",
x"A38C7CEA",
x"A2467C7C",
x"A0C07BE8",
x"9F0B7B22",
x"9D427A2C",
x"9B83790E",
x"99F377D7",
x"98B476A0",
x"97DA7583",
x"97777495",
x"978573E8",
x"97F67388",
x"98AB7375",
x"998173A7",
x"9A527410",
x"9AF6749C",
x"9B557534",
x"9B5F75CA",
x"9B14764B",
x"9A8576B0",
x"99CC76F8",
x"990A7722",
x"985F7731",
x"97E37729",
x"97A17706",
x"979076C6",
x"9795765A",
x"978175B7",
x"971874CB",
x"961E7388",
x"945771E2",
x"919D6FD8",
x"8DDD6D73",
x"89256AC5",
x"83A167EB",
x"7D9B650A",
x"77726249",
x"71895FD2",
x"6C455DC3",
x"67FA5C35",
x"64E35B2E",
x"63165AA9",
x"628C5A95",
x"631C5AD6",
x"64845B49",
x"667A5BCB",
x"68AE5C3D",
x"6AD95C90",
x"6CC55CB9",
x"6E525CBD",
x"6F775CAF",
x"70425CA4",
x"70CC5CB5",
x"71385CFD",
x"71AA5D8D",
x"72415E69",
x"730E5F91",
x"741E60F2",
x"75686274",
x"76DF63FD",
x"786D656C",
x"79FC66A7",
x"7B70679E",
x"7CBB6848",
x"7DCE68A4",
x"7EA168BB",
x"7F37689B",
x"7F936856",
x"7FBF6800",
x"7FC667A4",
x"7FB4674E",
x"7F906704",
x"7F6366C9",
x"7F32669A",
x"7F016675",
x"7ED16658",
x"7EA16641",
x"7E736630",
x"7E446627",
x"7E17662A",
x"7DEA663A",
x"7DC46656",
x"7DA46680",
x"7D9166B2",
x"7D9166EB",
x"7DA86720",
x"7DD9674C",
x"7E28676D",
x"7E93677C",
x"7F186777",
x"7FB26762",
x"8058673C",
x"80FA670D",
x"818E66D5",
x"8203669B",
x"82496660",
x"82586627",
x"822565ED",
x"81B265B2",
x"81016573",
x"8020652F",
x"7F1B64E2",
x"7E0D648D",
x"7D066431",
x"7C1D63D0",
x"7B5E6370",
x"7AD36314",
x"7A7C62C2",
x"7A526283",
x"7A49625A",
x"7A52624C",
x"7A5B625C",
x"7A566289",
x"7A3D62D2",
x"7A0D6331",
x"79C8639D",
x"797C640E",
x"7931647A",
x"78F764D5",
x"78D96515",
x"78DC6534",
x"78FF652B",
x"793B64FA",
x"798464A4",
x"79CC6431",
x"7A0263A7",
x"7A166311",
x"7A00627D",
x"79BB61F2",
x"79456179",
x"78A46114",
x"77E260C8",
x"77096090",
x"76246069",
x"753F604B",
x"74626032",
x"73936015",
x"72D65FF0",
x"72305FBF",
x"719D5F83",
x"711E5F3B",
x"70B05EE9",
x"70515E91",
x"6FFA5E39",
x"6FA85DE6",
x"6F555D9A",
x"6EFA5D59",
x"6E915D25",
x"6E165CFD",
x"6D845CE0",
x"6CDE5CCD",
x"6C205CBF",
x"6B535CB3",
x"6A7C5CA4",
x"69A05C8A",
x"68C75C63",
x"67F55C2B",
x"672B5BDD",
x"66695B77",
x"65AD5AFA",
x"64EF5A64",
x"642A59B9",
x"635758FD",
x"62705830",
x"6175575C",
x"60665684",
x"5F4A55B2",
x"5E2B54EB",
x"5D19543C",
x"5C2353AC",
x"5B5A5344",
x"5AD0530C",
x"5A8F5309",
x"5AA35340",
x"5B1053AD",
x"5BD15450",
x"5CDF551F",
x"5E2B5611",
x"5FA35718",
x"61335829",
x"62C45938",
x"64475A3C",
x"65AB5B2B",
x"66E95C02",
x"67FA5CC1",
x"68E35D64",
x"69AA5DEE",
x"6A565E60",
x"6AF55EBD",
x"6B905F07",
x"6C2E5F3F",
x"6CD45F67",
x"6D835F81",
x"6E355F92",
x"6EE65F9E",
x"6F8D5FA9",
x"701E5FB7",
x"70965FC8",
x"70ED5FDD",
x"71275FF9",
x"71486013",
x"7159602B",
x"7169603E",
x"71836048",
x"71B5604D",
x"720D6053",
x"72906060",
x"73416080",
x"741B60B8",
x"751A6113",
x"76316191",
x"77516232",
x"786C62ED",
x"797963B5",
x"7A6D647C",
x"7B476532",
x"7C0765CC",
x"7CB26642",
x"7D536696",
x"7DF266CB",
x"7E9666EF",
x"7F44670E",
x"7FFF6737",
x"80C16775",
x"818467C9",
x"823C6832",
x"82DE68A7",
x"835F6919",
x"83BB6977",
x"83F069B8",
x"840469D1",
x"840469C2",
x"84006994",
x"840B6958",
x"84396920",
x"849A6903",
x"85386916",
x"86146965",
x"872869F6",
x"88656AC2",
x"89B56BBE",
x"8AFE6CD4",
x"8C2A6DE9",
x"8D216EE9",
x"8DD66FC0",
x"8E42705F",
x"8E6770C1",
x"8E5270E9",
x"8E1070E2",
x"8DB470B9",
x"8D4F707A",
x"8CF07039",
x"8CA06FFC",
x"8C5C6FCA",
x"8C206FA0",
x"8BDF6F7C",
x"8B876F54",
x"8B0B6F1D",
x"8A5C6ECD",
x"89726E5B",
x"884B6DC1",
x"86ED6CFF",
x"85666C17",
x"83CC6B13",
x"823269FC",
x"80B268DE",
x"7F5F67C8",
x"7E4C66C5",
x"7D8165E2",
x"7D016525",
x"7CC96497",
x"7CCC6439",
x"7CF9640B",
x"7D3E6409",
x"7D86642F",
x"7DBF6477",
x"7DDB64DA",
x"7DD0654F",
x"7D9E65CE",
x"7D44664C",
x"7CC866C1",
x"7C34671E",
x"7B91675B",
x"7AE8676C",
x"7A3D6746",
x"799166E6",
x"78E06646",
x"7821656A",
x"774B6456",
x"7652631A",
x"752E61C3",
x"73D96067",
x"72565F18",
x"70AE5DE9",
x"6EF25CEC",
x"6D355C28",
x"6B945BA5",
x"6A275B61",
x"69095B56",
x"684B5B7A",
x"67F95BC0",
x"68165C1B",
x"689B5C81",
x"697D5CE9",
x"6AA75D4C",
x"6C045DA9",
x"6D7F5E03",
x"6F065E5A",
x"708A5EB7",
x"72045F1D",
x"73735F8E",
x"74D96011",
x"763B60A5",
x"779E614E",
x"790A620A",
x"7A8062D6",
x"7C0163B1",
x"7D876495",
x"7F0D6581",
x"8087666C",
x"81ED674F",
x"83356820",
x"845568D5",
x"85496966",
x"860D69CB",
x"86A16A02",
x"87076A09",
x"874369E3",
x"875C699D",
x"87556941",
x"873568E1",
x"87036889",
x"86C16849",
x"8671682B",
x"861A6831",
x"85BB685B",
x"8558689E",
x"84F368F3",
x"84936948",
x"843E6990",
x"83FD69C4",
x"83DC69DB",
x"83E669D5",
x"842569BC",
x"84A06999",
x"85566979",
x"8646696B",
x"87656979",
x"88A169AA",
x"89EA69FF",
x"8B2C6A75",
x"8C566B02",
x"8D596B9A",
x"8E2E6C31",
x"8ED56CB8",
x"8F526D26",
x"8FAF6D72",
x"8FF66D9A",
x"902C6D9D",
x"905C6D80",
x"90806D4A",
x"90956D02",
x"90946CB3",
x"906E6C65",
x"901E6C21",
x"8F9B6BED",
x"8EE66BD1",
x"8E046BCC",
x"8CFD6BE2",
x"8BE36C0F",
x"8AC46C4D",
x"89AE6C94",
x"88B16CDC",
x"87D56D1D",
x"871B6D4B",
x"86846D5E",
x"860D6D51",
x"85AC6D21",
x"855D6CD1",
x"85186C62",
x"84D56BDE",
x"848D6B49",
x"843C6AB0",
x"83DF6A13",
x"836F6979",
x"82E868E3",
x"82496851",
x"819067BB",
x"80BC6720",
x"7FD16679",
x"7ED265C6",
x"7DC86509",
x"7CBC6445",
x"7BBC6384",
x"7AD162D2",
x"7A04623E",
x"796361D3",
x"78F2619E",
x"78B461A4",
x"78AA61E6",
x"78D1625D",
x"791E62FD",
x"798663B2",
x"79F96469",
x"7A66650D",
x"7AB9658B",
x"7AE365D9",
x"7AD665F0",
x"7A8C65D0",
x"7A036584",
x"79416515",
x"78556495",
x"77516413",
x"76466395",
x"754B6328",
x"746862CB",
x"73A16276",
x"72F06221",
x"724561BF",
x"71866142",
x"7094609D",
x"6F515FC8",
x"6DA35EBC",
x"6B7A5D7B",
x"68D95C0E",
x"65CC5A7E",
x"627258DC",
x"5EF35738",
x"5B8355A5",
x"58555433",
x"559A52F7",
x"537951F8",
x"52095143",
x"515550DB",
x"515A50C4",
x"51FF50F7",
x"532B516E",
x"54B8521F",
x"568252FB",
x"586253F4",
x"5A3D54FA",
x"5BF955FF",
x"5D8856F8",
x"5EE257DA",
x"6007589C",
x"60FB593D",
x"61C559B9",
x"62735A14",
x"630F5A50",
x"63A35A76",
x"64375A8B",
x"64D25A9A",
x"65765AA6",
x"66275ABD",
x"66DF5AE3",
x"679B5B1A",
x"68555B63",
x"69035BBD",
x"699E5C1F",
x"6A215C82",
x"6A825CD9",
x"6ABD5D17",
x"6ACF5D31",
x"6ABA5D21",
x"6A805CE3",
x"6A265C7B",
x"69B45BF6",
x"69325B61",
x"68AD5AD2",
x"682B5A5C",
x"67BA5A12",
x"675F5A07",
x"67235A42",
x"67095AC5",
x"67135B87",
x"67415C7B",
x"67915D8E",
x"68005EA8",
x"688D5FB3",
x"6932609B",
x"69EF6152",
x"6AC161CE",
x"6BA4620D",
x"6C946211",
x"6D8D61E3",
x"6E86618E",
x"6F75611F",
x"704C60A2",
x"71006024",
x"71865FAC",
x"71D25F45",
x"71E25EF1",
x"71B45EB8",
x"714E5E9A",
x"70BA5E9A",
x"70095EB7",
x"6F4A5EED",
x"6E905F3F",
x"6DE95FA5",
x"6D63601D",
x"6D07609F",
x"6CD56124",
x"6CCC61A4",
x"6CE86218",
x"6D1E6279",
x"6D6662C1",
x"6DB562E9",
x"6E0462F2",
x"6E4C62D9",
x"6E8A62A2",
x"6EBA6250",
x"6EDC61E8",
x"6EF5616F",
x"6F0660ED",
x"6F13606A",
x"6F1D5FED",
x"6F255F78",
x"6F2D5F14",
x"6F2D5EBF",
x"6F215E7A",
x"6F025E45",
x"6EC55E1A",
x"6E665DF7",
x"6DDF5DD5",
x"6D2E5DB2",
x"6C595D87",
x"6B695D53",
x"6A6D5D12",
x"697B5CC8",
x"68A35C71",
x"67FC5C14",
x"67915BB2",
x"67705B52",
x"67945AFA",
x"67F85AAE",
x"68895A76",
x"69305A56",
x"69D65A4F",
x"6A625A60",
x"6ABE5A88",
x"6ADB5ABD",
x"6AB05AF8",
x"6A3F5B2C",
x"69915B4D",
x"68B55B52",
x"67BE5B33",
x"66C15AF0",
x"65D15A8B",
x"64FC5A0B",
x"644E5980",
x"63CB58F7",
x"636F5880",
x"63305825",
x"62FF57ED",
x"62CB57D7",
x"628057DC",
x"620D57EE",
x"616557FE",
x"607F57FA",
x"5F5E57D1",
x"5E0C577F",
x"5C9A5702",
x"5B235660",
x"59C755A8",
x"58A454EE",
x"57D95449",
x"577F53CA",
x"57A15382",
x"5844537D",
x"595E53B6",
x"5ADA542D",
x"5C9A54D3",
x"5E7D5599",
x"605E5671",
x"621A574A",
x"639A581C",
x"64C858E0",
x"65A15995",
x"66245A3D",
x"665E5ADF",
x"665E5B7D",
x"66385C1A",
x"66035CB8",
x"65CE5D50",
x"65A75DDF",
x"65965E55",
x"65A05EAB",
x"65C45ED6",
x"66025ECF",
x"66545E94",
x"66B75E28",
x"672D5D95",
x"67B35CE9",
x"68485C35",
x"68ED5B8E",
x"69A15B04",
x"6A5C5AA8",
x"6B195A81",
x"6BCB5A92",
x"6C665ADA",
x"6CDE5B4C",
x"6D275BD9",
x"6D385C71",
x"6D115D01",
x"6CB45D7B",
x"6C2A5DD2",
x"6B825E00",
x"6ACC5E04",
x"6A1C5DE3",
x"69825DA7",
x"69075D5A",
x"68B45D0B",
x"68895CC5",
x"687F5C91",
x"688D5C73",
x"68A85C6E",
x"68CA5C81",
x"68E85CA4",
x"69025CD2",
x"69195D02",
x"69345D2F",
x"695C5D52",
x"69995D67",
x"69F05D70",
x"6A635D6E",
x"6AED5D69",
x"6B845D62",
x"6C1D5D5F",
x"6CA35D63",
x"6D075D71",
x"6D3E5D86",
x"6D3B5D9B",
x"6CFD5DA9",
x"6C8C5DA8",
x"6BEF5D8E",
x"6B3A5D56",
x"6A7F5D00",
x"69CF5C8E",
x"69415C0B",
x"68DE5B85",
x"68B05B0E",
x"68B75AB6",
x"68F25A90",
x"69585AA4",
x"69DF5AFA",
x"6A7A5B8E",
x"6B1E5C57",
x"6BC15D48",
x"6C585E4B",
x"6CDE5F4C",
x"6D516038",
x"6DAE6100",
x"6DF86197",
x"6E2D61F3",
x"6E516215",
x"6E6561FD",
x"6E6961AF",
x"6E5F6131",
x"6E45608A",
x"6E1B5FC5",
x"6DDF5EE7",
x"6D905DFE",
x"6D2D5D14",
x"6CB35C32",
x"6C215B66",
x"6B795AB6",
x"6AB85A2F",
x"69E159D2",
x"68F5599E",
x"67F95992",
x"66F659A5",
x"65F659CC",
x"650259FB",
x"642A5A26",
x"63795A45",
x"62FB5A53",
x"62B75A4F",
x"62AE5A3D",
x"62DE5A25",
x"63385A0E",
x"63AA59FE",
x"641959F8",
x"646659FB",
x"64795A01",
x"64345A00",
x"638659EA",
x"626859B0",
x"60DE594A",
x"5EFA58B3",
x"5CDB57EB",
x"5AA756FF",
x"588C5602",
x"56B8550F",
x"55525440",
x"547C53B2",
x"544A537A",
x"54C153A5",
x"55D55433",
x"5773551B",
x"59765644",
x"5BBA5791",
x"5E1258DD",
x"60565A07",
x"62695AF0",
x"64315B87",
x"65A05BC6",
x"66B45BB6",
x"67755B6A",
x"67F25B00",
x"683D5A97",
x"686C5A4F",
x"68905A3D",
x"68BB5A70",
x"68F55AE9",
x"69415B9A",
x"699C5C6E",
x"69FF5D4C",
x"6A5B5E15",
x"6AA75EB3",
x"6AD85F15",
x"6AE65F37",
x"6AD45F1D",
x"6AA35ED6",
x"6A5F5E7A",
x"6A1A5E1E",
x"69E65DD9",
x"69D55DB6",
x"69F35DBD",
x"6A485DED",
x"6AD45E39",
x"6B8D5E95",
x"6C655EED",
x"6D445F35",
x"6E135F63",
x"6EBB5F74",
x"6F2E5F6D",
x"6F635F59",
x"6F5E5F45",
x"6F275F3F",
x"6ED45F53",
x"6E7C5F8A",
x"6E3A5FE2",
x"6E206053",
x"6E3E60D3",
x"6E9A6152",
x"6F2E61BF",
x"6FED620B",
x"70C8622F",
x"71A76228",
x"727961F9",
x"733261AD",
x"73CE6155",
x"744F6104",
x"74BE60CC",
x"752A60BE",
x"759E60E4",
x"76256142",
x"76C661D5",
x"777C6294",
x"783C6370",
x"78F66456",
x"79966534",
x"7A0765F7",
x"7A3B6690",
x"7A2766F6",
x"79CC6723",
x"79316716",
x"786566D8",
x"777D666F",
x"768F65E8",
x"75AE654C",
x"74EC64AA",
x"7452640B",
x"73E66376",
x"73A462F3",
x"73876284",
x"7387622E",
x"739A61EF",
x"73B761C8",
x"73D961B5",
x"73FC61B5",
x"741E61C2",
x"743D61D6",
x"745B61EA",
x"747361F6",
x"748661F3",
x"748E61DA",
x"748761A7",
x"746C6155",
x"743760E7",
x"73E66063",
x"73785FCF",
x"72EC5F35",
x"72475E9F",
x"718C5E1C",
x"70C15DB5",
x"6FEF5D70",
x"6F1B5D53",
x"6E4F5D5A",
x"6D915D84",
x"6CE95DC6",
x"6C595E15",
x"6BE65E66",
x"6B935EAB",
x"6B5B5ED9",
x"6B385EEA",
x"6B245ED7",
x"6B105EA2",
x"6AED5E4C",
x"6AAB5DD6",
x"6A3B5D48",
x"698D5CA4",
x"68975BEE",
x"67565B29",
x"65CB5A57",
x"63FD597A",
x"61FF588F",
x"5FE1579C",
x"5DC056A5",
x"5BB755B0",
x"59E254C7",
x"585E53F4",
x"57415343",
x"569D52BF",
x"567C5271",
x"56E25263",
x"57CA5295",
x"59235309",
x"5ADB53BC",
x"5CD754A6",
x"5EFA55BF",
x"612A56FB",
x"634B5850",
x"654859B2",
x"67145B15",
x"68A85C6D",
x"6A055DB1",
x"6B315ED7",
x"6C3B5FD9",
x"6D3360B4",
x"6E276163",
x"6F2461EC",
x"70346252",
x"7155629D",
x"728762D2",
x"73BE62FC",
x"74EC631F",
x"76036342",
x"76F56362",
x"77B5637F",
x"783E6395",
x"789063A3",
x"78B163A1",
x"78AA6393",
x"788A6379",
x"78626359",
x"783C633E",
x"7826632B",
x"7822632D",
x"78306344",
x"784B6373",
x"786963B8",
x"7880640B",
x"78896462",
x"787C64B5",
x"785B64FC",
x"782A6531",
x"77F66553",
x"77CE6566",
x"77C16572",
x"77DD657A",
x"782D6589",
x"78B065A3",
x"796365C8",
x"7A3865F7",
x"7B1E662E",
x"7BFD6660",
x"7CBF668A",
x"7D5066A4",
x"7DA566A8",
x"7DB56699",
x"7D846676",
x"7D1B6646",
x"7C8B6613",
x"7BE565E3",
x"7B3C65BF",
x"7AA365AD",
x"7A2165AF",
x"79C265C8",
x"798465F3",
x"7968662E",
x"79636673",
x"797266BA",
x"798C66FC",
x"79A86731",
x"79C76753",
x"79E3675C",
x"79FF674B",
x"7A18671A",
x"7A3166CE",
x"7A496669",
x"7A5D65F5",
x"7A6C6579",
x"7A706500",
x"7A666497",
x"7A496448",
x"7A18641A",
x"79D26411",
x"7977642A",
x"790C645F",
x"789164A7",
x"780E64F2",
x"77846534",
x"76F9655E",
x"766C6568",
x"75E06549",
x"75556503",
x"74CF6498",
x"744E6414",
x"73D86380",
x"737262EC",
x"73216264",
x"72ED61FA",
x"72DC61B1",
x"72F26191",
x"732E6198",
x"738E61C2",
x"740D6206",
x"74A06258",
x"753A62AB",
x"75CE62F4",
x"764F632A",
x"76B26346",
x"76EC6346",
x"76F9632E",
x"76D56301",
x"768062C5",
x"75FD6281",
x"754F623B",
x"747C61F4",
x"738461A9",
x"726F6158",
x"713A60F6",
x"6FE9607C",
x"6E7C5FE2",
x"6CF55F22",
x"6B535E3D",
x"69A05D39",
x"67DE5C1C",
x"66195AF6",
x"645E59D3",
x"62BB58C6",
x"614457DC",
x"6009571E",
x"5F1A5694",
x"5E88563D",
x"5E595618",
x"5E93561C",
x"5F335642",
x"602B5681",
x"616E56D0",
x"62E3572C",
x"6476578F",
x"660C57F8",
x"678F5869",
x"68EF58E1",
x"6A205964",
x"6B1E59F1",
x"6BEF5A88",
x"6C9A5B29",
x"6D2B5BD3",
x"6DB35C84",
x"6E3B5D39",
x"6ECF5DF1",
x"6F755EAC",
x"702D5F6C",
x"70F3602D",
x"71C160F2",
x"728D61B8",
x"734F6280",
x"74006345",
x"749B6403",
x"751E64B2",
x"758C654C",
x"75E365C9",
x"762E6623",
x"76706653",
x"76B06659",
x"76F26638",
x"773865F2",
x"77876591",
x"77DF6521",
x"783C64AD",
x"78A16441",
x"790763E5",
x"797063A1",
x"79D86379",
x"7A3E636D",
x"7AA4637A",
x"7B0A639B",
x"7B7363CE",
x"7BE5640A",
x"7C5F6450",
x"7CE5649D",
x"7D7964F3",
x"7E176553",
x"7EBC65BF",
x"7F63663A",
x"800166C1",
x"80906755",
x"810667F0",
x"8160688E",
x"819E692A",
x"81C269BE",
x"81D56A44",
x"81E26ABA",
x"81F96B1E",
x"82256B72",
x"82746BB5",
x"82EC6BEC",
x"838A6C13",
x"84466C2D",
x"85116C35",
x"85D36C2D",
x"86736C0F",
x"86D86BDB",
x"86EC6B8D",
x"86A16B2A",
x"85F36AB1",
x"84E76A28",
x"838E6996",
x"820368FD",
x"80626866",
x"7ECC67D8",
x"7D5F6753",
x"7C3266DE",
x"7B536676",
x"7AC56620",
x"7A8265D8",
x"7A77659E",
x"7A8E6572",
x"7AAE654F",
x"7ABB6535",
x"7AA16523",
x"7A536513",
x"79CC6501",
x"791164ED",
x"783164D2",
x"773F64AE",
x"76566483",
x"758F6450",
x"74FF641A",
x"74B763E0",
x"74BE63AB",
x"7513637A",
x"75A56352",
x"76656331",
x"77356318",
x"77FC6304",
x"789B62F4",
x"790162E3",
x"792062CF",
x"78F562B7",
x"78846298",
x"77DF6274",
x"7717624B",
x"7644621B",
x"757661E2",
x"74B8619B",
x"740C6141",
x"736960CB",
x"72BE6033",
x"71F35F74",
x"70F25E8A",
x"6FA35D7A",
x"6DFD5C48",
x"6C005B01",
x"69BB59B8",
x"674B587D",
x"64D45764",
x"62855681",
x"608755E1",
x"5F04558C",
x"5E175584",
x"5DCE55C6",
x"5E295649",
x"5F1C5701",
x"608D57E0",
x"626258D7",
x"647959DC",
x"66B75AE3",
x"69025BE9",
x"6B4B5CE9",
x"6D845DE2",
x"6FA85ED5",
x"71B55FC1",
x"73A860A5",
x"757F6181",
x"77376255",
x"78CB631D",
x"7A3863D8",
x"7B7A6483",
x"7C936520",
x"7D8465B1",
x"7E536638",
x"7F0966BA",
x"7FB16738",
x"805267B7",
x"80F66834",
x"81A068B0",
x"82506926",
x"83036994",
x"83AF69F6",
x"844F6A45",
x"84D66A83",
x"853C6AAE",
x"857F6AC8",
x"859B6AD5",
x"85956AD9",
x"85766ADC",
x"85446AE2",
x"850B6AF0",
x"84DA6B07",
x"84B86B2D",
x"84B16B5F",
x"84C66B9E",
x"85006BEB",
x"855B6C44",
x"85D36CAA",
x"86676D1D",
x"870E6DA0",
x"87BF6E30",
x"88726ECE",
x"891A6F78",
x"89AE7027",
x"8A2570D7",
x"8A76717E",
x"8A9D7213",
x"8A9A728C",
x"8A7072E1",
x"8A297309",
x"89D57303",
x"898172D2",
x"89417279",
x"89247205",
x"89387183",
x"89817105",
x"8A037096",
x"8AAF7047",
x"8B76701A",
x"8C407014",
x"8CF6702E",
x"8D7A705A",
x"8DBB7088",
x"8DAA70A4",
x"8D4270A1",
x"8C8D7073",
x"8B987013",
x"8A7E6F88",
x"89586EDB",
x"88416E20",
x"87526D6E",
x"869B6CD7",
x"86256C6F",
x"85ED6C3E",
x"85EC6C47",
x"86116C80",
x"864C6CDF",
x"868B6D4E",
x"86C16DBA",
x"86E66E10",
x"86F76E44",
x"86FA6E52",
x"86F76E38",
x"86FC6E00",
x"87126DB5",
x"87456D63",
x"87976D19",
x"880A6CDB",
x"88986CB3",
x"89386C9D",
x"89DC6C9A",
x"8A776CA3",
x"8AFB6CB1",
x"8B626CC1",
x"8BA16CCF",
x"8BB66CDE",
x"8BA16CEE",
x"8B676D00",
x"8B106D1A",
x"8AA26D3B",
x"8A2B6D65",
x"89B16D93",
x"893F6DC1",
x"88DA6DE6",
x"88866DFD",
x"88416DFC",
x"88006DD9",
x"87B56D8F",
x"874B6D16",
x"86A56C69",
x"85A56B82",
x"842E6A5C",
x"822368F7",
x"7F736752",
x"7C1B6570",
x"78266359",
x"73AB6118",
x"6ED85EC1",
x"69E25C67",
x"65085A26",
x"60895815",
x"5C9E564D",
x"597B54E1",
x"573D53DD",
x"55F15343",
x"55925311",
x"56095339",
x"573053AB",
x"58DA5453",
x"5AD1551B",
x"5CE955F3",
x"5EF356CF",
x"60D257A8",
x"626F587E",
x"63C25953",
x"64CF5A2E",
x"65A45B12",
x"66555C06",
x"66FC5D0A",
x"67B15E1A",
x"688A5F32",
x"69996048",
x"6AE26152",
x"6C666246",
x"6E19631D",
x"6FE663CE",
x"71B76456",
x"737264B7",
x"74FC64F2",
x"7645650D",
x"773E650D",
x"77E864FD",
x"784664E3",
x"786964C9",
x"786564B7",
x"784E64AF",
x"783864B7",
x"783464CE",
x"784964F4",
x"78796528",
x"78BF6566",
x"791465A8",
x"796C65ED",
x"79BE6635",
x"7A066681",
x"7A4566D3",
x"7A836731",
x"7AC7679A",
x"7B1E6811",
x"7B986893",
x"7C3C6917",
x"7D106996",
x"7E106A02",
x"7F346A4F",
x"806C6A73",
x"81A76A6B",
x"82CF6A37",
x"83D269E2",
x"84A16979",
x"852F6911",
x"857B68BC",
x"8589688A",
x"855C6884",
x"850368AB",
x"848968F7",
x"83FC6956",
x"836969B5",
x"82D969FF",
x"82526A1D",
x"81D96A09",
x"817269BC",
x"81186941",
x"80D168A4",
x"809767FF",
x"806F6763",
x"805666E5",
x"804F6693",
x"8059666F",
x"80736675",
x"809B669A",
x"80CB66CC",
x"80FA66FC",
x"81226717",
x"81386714",
x"813166F0",
x"810366AD",
x"80A76650",
x"801A65E6",
x"7F5C6579",
x"7E726513",
x"7D5F64B7",
x"7C326468",
x"7AF66421",
x"79B763DF",
x"7884639D",
x"776B6353",
x"76756304",
x"75B162B1",
x"7524625F",
x"74D66217",
x"74C961E3",
x"74FF61CE",
x"756F61DC",
x"76146214",
x"76E26272",
x"77C662F3",
x"78B4638D",
x"79966439",
x"7A5D64EA",
x"7AFE6597",
x"7B726638",
x"7BB566C9",
x"7BCC6744",
x"7BBF67A8",
x"7B9767F5",
x"7B5E6826",
x"7B18683C",
x"7AC86831",
x"7A666801",
x"79E667A5",
x"79346717",
x"78386652",
x"76E06552",
x"7517641A",
x"72D562AE",
x"701B6114",
x"6CF95F5A",
x"69875D8E",
x"65EB5BBF",
x"624F5A00",
x"5EE5585D",
x"5BD756E6",
x"594A55A6",
x"575954A3",
x"561453E7",
x"557B5370",
x"5580533D",
x"560F534E",
x"570A539C",
x"5851541F",
x"59C554CA",
x"5B4A5591",
x"5CCB5666",
x"5E3A5739",
x"5F8F57FD",
x"60C758A6",
x"61E6592E",
x"62F1598F",
x"63EB59D2",
x"64DB59FE",
x"65BF5A21",
x"669B5A4D",
x"676B5A92",
x"682B5AFE",
x"68D85B9B",
x"696B5C69",
x"69E15D5F",
x"6A385E70",
x"6A6D5F86",
x"6A826087",
x"6A75615F",
x"6A4B61F7",
x"6A076245",
x"69B16243",
x"694F61FA",
x"68E86176",
x"688760CE",
x"6833601B",
x"67F55F74",
x"67D25EF3",
x"67D15EA4",
x"67F05E90",
x"68335EB8",
x"68915F12",
x"69075F95",
x"698F602E",
x"6A2160CE",
x"6AB86160",
x"6B5261DD",
x"6BEF623B",
x"6C906277",
x"6D3A6291",
x"6DF3628E",
x"6EBF6274",
x"6F9E624C",
x"7090621A",
x"718D61E6",
x"728A61B5",
x"73766188",
x"74426164",
x"74DE614B",
x"753A6139",
x"75516132",
x"75206138",
x"74B26148",
x"74166163",
x"73636188",
x"72B161B8",
x"721D61EF",
x"71BE622B",
x"71A4626A",
x"71D862A8",
x"725962E3",
x"731D631A",
x"740E6349",
x"75166372",
x"761A6393",
x"770163AD",
x"77B863C1",
x"783163CF",
x"786563D6",
x"785963D6",
x"781763CF",
x"77B263BC",
x"773E639E",
x"76CB6370",
x"766F6332",
x"763562E6",
x"7624628A",
x"763F6222",
x"767F61B4",
x"76DB6145",
x"774560DC",
x"77B2607E",
x"78136037",
x"785C6007",
x"78895FF6",
x"78986003",
x"788A602E",
x"78676076",
x"783A60D5",
x"78076142",
x"77DB61B5",
x"77BA6225",
x"77A56287",
x"779A62D2",
x"779462FD",
x"778A6304",
x"777562EA",
x"774C62AF",
x"770E625F",
x"76BA6203",
x"765461A8",
x"75DF615D",
x"75636129",
x"74E26113",
x"74586113",
x"73BE6122",
x"7304612F",
x"721C6125",
x"70F360EE",
x"6F7F6079",
x"6DBE5FBB",
x"6BBD5EB8",
x"69995D7B",
x"677A5C22",
x"659C5AD0",
x"643559B0",
x"638258EA",
x"63AE58A4",
x"64D758F3",
x"670059E1",
x"6A165B69",
x"6DEE5D71",
x"724B5FDA",
x"76E86277",
x"7B7D6520",
x"7FCB67A7",
x"83A169F0",
x"86E06BE2",
x"897D6D75",
x"8B816EA7",
x"8D066F85",
x"8E28701C",
x"8F107082",
x"8FE370CE",
x"90C27116",
x"91C9716E",
x"930E71E6",
x"949B7292",
x"967A7379",
x"98A874A3",
x"9B21760C",
x"9DD677AF",
x"A0B6797C",
x"A3A67B60",
x"A68D7D3F",
x"A9497EFF",
x"ABBC808B",
x"ADCF81CD",
x"AF7182B8",
x"B09C834A",
x"B156838E",
x"B1AF8392",
x"B1C28370",
x"B1AB8342",
x"B18B831F",
x"B17E831C",
x"B1988345",
x"B1E18399",
x"B25D8415",
x"B30184A8",
x"B3C38543",
x"B48F85D6",
x"B5598650",
x"B61486AB",
x"B6BA86E6",
x"B74C8705",
x"B7CD8715",
x"B8498725",
x"B8C78743",
x"B953877D",
x"B9F487D9",
x"BAAD8859",
x"BB7D88F9",
x"BC5B89A9",
x"BD3C8A5D",
x"BE0F8B00",
x"BEC18B7D",
x"BF3F8BC8",
x"BF748BD2",
x"BF4F8B97",
x"BEC78B18",
x"BDD98A5F",
x"BC888977",
x"BAE68873",
x"B90A8766",
x"B7158660",
x"B5298577",
x"B36E84B9",
x"B2078431",
x"B10A83E8",
x"B08A83E1",
x"B088841B",
x"B0FD848F",
x"B1CF8535",
x"B2DE85FD",
x"B40786D9",
x"B52287B3",
x"B609887D",
x"B6A28922",
x"B6D98995",
x"B6A589CC",
x"B60C89BF",
x"B51B8970",
x"B3E188E2",
x"B2778819",
x"B0F08725",
x"AF60860D",
x"ADD384DC",
x"AC528399",
x"AAD9824D",
x"A9698100",
x"A7FB7FB5",
x"A68B7E72",
x"A5147D3C",
x"A3987C1B",
x"A21C7B15",
x"A0A97A33",
x"9F4A7978",
x"9E0A78E7",
x"9CF7787F",
x"9C17783C",
x"9B6E7812",
x"9AFD77F8",
x"9AB877E1",
x"9A9777C3",
x"9A8A7796",
x"9A837757",
x"9A77770C",
x"9A6076BC",
x"9A3C7678",
x"9A14764E",
x"99F07652",
x"99DC768F",
x"99E7770D",
x"9A1777CA",
x"9A6B78BA",
x"9AD979C7",
x"9B467AD3",
x"9B917BB7",
x"9B8E7C4C",
x"9B0E7C68",
x"99E77BEF",
x"97F67AC9",
x"952978ED",
x"91857661",
x"8D247340",
x"88376FAE",
x"82FD6BDF",
x"7DC5680A",
x"78DC6469",
x"748C612F",
x"710D5E8A",
x"6E845C94",
x"6D005B5C",
x"6C795ADF",
x"6CD45B0D",
x"6DE85BCB",
x"6F8A5CFA",
x"718E5E77",
x"73CC6024",
x"762861E3",
x"789063A4",
x"7AF76556",
x"7D5C66F6",
x"7FBA687C",
x"820E69E8",
x"84566B3A",
x"86866C72",
x"88916D8C",
x"8A6F6E86",
x"8C136F5F",
x"8D797013",
x"8EA270A4",
x"8F947114",
x"905C7166",
x"910671A3",
x"91A171CF",
x"923C71F4",
x"92DF7216",
x"938B723B",
x"94437266",
x"94FE7297",
x"95B572D0",
x"9660730B",
x"96F67347",
x"97707380",
x"97CD73B4",
x"980B73DE",
x"982873FB",
x"98257406",
x"980473FF",
x"97C573E1",
x"976A73AA",
x"96F8735E",
x"967672FB",
x"95EA7288",
x"9563720C",
x"94EF718F",
x"949F711D",
x"948770C3",
x"94B97089",
x"95437078",
x"962F7097",
x"977E70E9",
x"992B716B",
x"9B257215",
x"9D5372E1",
x"9F9873C3",
x"A1D074AD",
x"A3D77593",
x"A58D766C",
x"A6D6772C",
x"A79C77CB",
x"A7DC7844",
x"A7957892",
x"A6DA78B6",
x"A5BF78B0",
x"A4647882",
x"A2EB7834",
x"A17377CD",
x"A0177752",
x"9EEC76D1",
x"9DFD7652",
x"9D4D75DC",
x"9CD77578",
x"9C8B752A",
x"9C5C74F5",
x"9C3574DA",
x"9C0A74D4",
x"9BCB74E5",
x"9B717506",
x"9AFA7534",
x"9A64756E",
x"99B475AF",
x"98E975F4",
x"980D763A",
x"9721767B",
x"962976B1",
x"952976D4",
x"942576D8",
x"932176B4",
x"921E7660",
x"912475D4",
x"90357510",
x"8F537416",
x"8E8372F1",
x"8DC271AF",
x"8D0D7061",
x"8C626F1D",
x"8BB86DF8",
x"8B106D02",
x"8A646C48",
x"89B56BCF",
x"89046B96",
x"88566B90",
x"87B16BB1",
x"87166BE2",
x"86886C12",
x"86066C27",
x"858A6C13",
x"850A6BCB",
x"847C6B49",
x"83D36A90",
x"830669A6",
x"820D6899",
x"80E56779",
x"7F8D6656",
x"7E0B653F",
x"7C66643E",
x"7AA36356",
x"78C5628A",
x"76CC61CF",
x"74B8611F",
x"7282606C",
x"70245FAB",
x"6D9B5ED2",
x"6AEB5DDC",
x"681B5CCD",
x"65415BAE",
x"62785A8A",
x"5FE25974",
x"5DA75880",
x"5BE957C2",
x"5ACB5747",
x"5A5E571C",
x"5AAA573F",
x"5BA957AC",
x"5D425856",
x"5F55592C",
x"61B85A1B",
x"64415B0E",
x"66C45BF3",
x"69205CBD",
x"6B3E5D66",
x"6D165DEC",
x"6EA45E55",
x"6FF65EA9",
x"711B5EF7",
x"72285F49",
x"732E5FAB",
x"743F6025",
x"756260BC",
x"769B6172",
x"77E56242",
x"79356327",
x"7A806417",
x"7BB96509",
x"7CD465F5",
x"7DC566D2",
x"7E896797",
x"7F216842",
x"7F9068CF",
x"7FE2693E",
x"80216990",
x"805969C9",
x"809A69F0",
x"80ED6A0A",
x"81566A1D",
x"81D66A2D",
x"82696A41",
x"83046A5C",
x"83986A7D",
x"84116AA6",
x"84606AD2",
x"84766AFD",
x"84486B24",
x"83D86B44",
x"832E6B57",
x"825A6B5C",
x"81776B58",
x"809E6B4B",
x"7FEF6B3A",
x"7F806B2D",
x"7F636B28",
x"7F9D6B32",
x"80276B4E",
x"80EF6B7C",
x"81D86BBA",
x"82C46C02",
x"838E6C4D",
x"841B6C8D",
x"84566CBB",
x"84376CCB",
x"83BF6CB4",
x"83006C72",
x"82106C03",
x"810E6B6F",
x"80186ABD",
x"7F4969FA",
x"7EBA693B",
x"7E736890",
x"7E7C680E",
x"7ECE67C5",
x"7F5D67BF",
x"801A6804",
x"80F26893",
x"81D56961",
x"82B26A5E",
x"83836B78",
x"843E6C92",
x"84E06D96",
x"85696E69",
x"85DC6EFC",
x"86366F3E",
x"867D6F2E",
x"86AB6ED1",
x"86C16E31",
x"86BB6D62",
x"86986C7A",
x"86566B94",
x"85F76AC2",
x"857F6A17",
x"84EF699D",
x"84506956",
x"83AE6941",
x"83106952",
x"827D697D",
x"820169B2",
x"819E69E5",
x"815B6A0A",
x"81356A1E",
x"812D6A1D",
x"813B6A0A",
x"815D69EC",
x"818869C7",
x"81B869A1",
x"81E0697F",
x"81FC695F",
x"82036942",
x"81F06924",
x"81BE6900",
x"816A68D1",
x"80F66894",
x"805F6849",
x"7FA867ED",
x"7ED26783",
x"7DDD670B",
x"7CCC6686",
x"7B9D65F5",
x"7A4E6552",
x"78E0649E",
x"775563D6",
x"75AE62F9",
x"73F26207",
x"72306106",
x"70766000",
x"6EDC5F00",
x"6D7D5E1A",
x"6C755D5D",
x"6BDC5CDD",
x"6BCC5CA8",
x"6C535CC9",
x"6D795D43",
x"6F3A5E15",
x"71865F37",
x"7448609B",
x"7763622F",
x"7AB863E3",
x"7E2465A3",
x"818B675E",
x"84D86907",
x"87F96A97",
x"8AE76C0A",
x"8DA86D62",
x"90426EA4",
x"92C56FD9",
x"9542710C",
x"97C9724A",
x"9A69739C",
x"9D2B750C",
x"A00F76A0",
x"A3117856",
x"A6217A26",
x"A9267C06",
x"AC077DE0",
x"AE9E7F9E",
x"B0CF8126",
x"B27A8266",
x"B3888347",
x"B3F183C2",
x"B3B683D7",
x"B2E68391",
x"B19F8304",
x"B007824C",
x"AE4C818A",
x"ACA180DB",
x"AB2D805D",
x"AA1C8022",
x"A9858033",
x"A97D808F",
x"AA05812C",
x"AB1981FD",
x"ACAD82EB",
x"AEAE83EA",
x"B10884EC",
x"B3A385EC",
x"B66A86EA",
x"B94387EE",
x"BC198901",
x"BED38A29",
x"C1588B6D",
x"C3938CC8",
x"C5718E32",
x"C6E08F9E",
x"C7DB90F7",
x"C865922B",
x"C88E9327",
x"C86A93DC",
x"C8189448",
x"C7BD946C",
x"C77B9452",
x"C770940A",
x"C7AF93A7",
x"C843933B",
x"C92592D6",
x"CA4A9287",
x"CB999252",
x"CCF59238",
x"CE439237",
x"CF679245",
x"D04B9258",
x"D0E59266",
x"D12D9265",
x"D126924C",
x"D0D79216",
x"D04A91C1",
x"CF8F9151",
x"CEB790C9",
x"CDD79037",
x"CD018FA8",
x"CC498F2F",
x"CBC18EDC",
x"CB7B8EC1",
x"CB818EE9",
x"CBD58F5B",
x"CC759016",
x"CD519110",
x"CE549238",
x"CF619378",
x"D05A94B1",
x"D12095CC",
x"D19C96B0",
x"D1C3974B",
x"D1929797",
x"D1199796",
x"D071974E",
x"CFB996D4",
x"CF199638",
x"CEB19590",
x"CE9B94EF",
x"CEE2945F",
x"CF8893EA",
x"D0779390",
x"D192934C",
x"D2B09311",
x"D3A592D6",
x"D443928C",
x"D4619223",
x"D3E49190",
x"D2B790C8",
x"D0D88FC6",
x"CE508E89",
x"CB338D0D",
x"C79D8B5C",
x"C3B0897B",
x"BF898776",
x"BB438559",
x"B6F1832C",
x"B29880FB",
x"AE307EC9",
x"A9AB7C91",
x"A4E97A4B",
x"9FC977EE",
x"9A317568",
x"940872AA",
x"8D4D6FA7",
x"860D6C5F",
x"7E6D68D8",
x"76AB6524",
x"6F166162",
x"68055DBB",
x"61D25A5A",
x"5CD2576E",
x"5940551C",
x"57405382",
x"56D552AF",
x"57E852A5",
x"5A3D5354",
x"5D8A54A5",
x"617B5675",
x"65B5589E",
x"69ED5AF8",
x"6DE35D64",
x"71725FC2",
x"748361FC",
x"771A63FF",
x"794765C4",
x"7B236744",
x"7CC86880",
x"7E53697A",
x"7FD86A3B",
x"815D6ACC",
x"82E66B3B",
x"846C6B97",
x"85E36BEF",
x"873C6C52",
x"886F6CCA",
x"896F6D5C",
x"8A376E09",
x"8AC96ECA",
x"8B2E6F93",
x"8B6C7055",
x"8B947100",
x"8BB17183",
x"8BCF71D2",
x"8BF771E8",
x"8C3271C1",
x"8C7E7164",
x"8CDA70DA",
x"8D3F7030",
x"8DA56F75",
x"8E006EB8",
x"8E486E06",
x"8E776D6B",
x"8E876CEC",
x"8E796C92",
x"8E4F6C5C",
x"8E116C4E",
x"8DC66C63",
x"8D776C99",
x"8D2B6CE6",
x"8CE96D45",
x"8CB46DA9",
x"8C8D6E06",
x"8C706E54",
x"8C5A6E89",
x"8C4B6EA4",
x"8C3C6EA4",
x"8C2F6E8D",
x"8C256E69",
x"8C216E44",
x"8C286E27",
x"8C426E20",
x"8C736E35",
x"8CC26E6C",
x"8D316EC4",
x"8DBF6F38",
x"8E6A6FC4",
x"8F2C705C",
x"900070FE",
x"90DA71A0",
x"91B57240",
x"928872DE",
x"934C737B",
x"93FB7416",
x"949174AF",
x"950B7546",
x"956975D5",
x"95AC7657",
x"95D576C3",
x"95E97710",
x"95E97737",
x"95DA7731",
x"95C276FE",
x"95A476A0",
x"9588761F",
x"95717586",
x"956974E5",
x"9574744D",
x"959873CB",
x"95DF7372",
x"964B734E",
x"96E27368",
x"97A273C3",
x"988A745E",
x"99927537",
x"9AAF7641",
x"9BD0776F",
x"9CE778B0",
x"9DE279EF",
x"9EB17B1C",
x"9F497C20",
x"9FA57CED",
x"9FC57D72",
x"9FAB7DA9",
x"9F637D8F",
x"9EF77D25",
x"9E747C71",
x"9DE67B85",
x"9D567A6E",
x"9CCC7943",
x"9C4F7816",
x"9BE376FE",
x"9B907609",
x"9B597548",
x"9B4074C1",
x"9B4B7476",
x"9B737462",
x"9BAF7479",
x"9BEE74A7",
x"9C1174D7",
x"9BF674EB",
x"9B7074CA",
x"9A567458",
x"98837380",
x"95DA7234",
x"92587070",
x"8E046E3A",
x"89046BA4",
x"839168CE",
x"7DF365DB",
x"787C62F7",
x"737F6052",
x"6F475E14",
x"6C0E5C60",
x"69FC5B50",
x"691E5AEE",
x"69685B38",
x"6ABB5C1E",
x"6CE65D84",
x"6FB05F4B",
x"72DF614C",
x"763B6366",
x"79976576",
x"7CD06766",
x"7FD36926",
x"82976AAE",
x"851A6C00",
x"87636D23",
x"897C6E23",
x"8B6A6F0C",
x"8D346FEC",
x"8EDC70CE",
x"906371BB",
x"91C572B7",
x"92FD73C0",
x"940A74D2",
x"94E775E5",
x"959776EB",
x"961777D7",
x"9669789B",
x"96907925",
x"968A796B",
x"96557964",
x"95F0790E",
x"9556786A",
x"94867781",
x"937E7662",
x"92487525",
x"90EA73DB",
x"8F7A729F",
x"8E0B7188",
x"8CBB70A6",
x"8BA27008",
x"8ADC6FB3",
x"8A7D6FA4",
x"8A906FD5",
x"8B177035",
x"8C0B70B3",
x"8D5D713B",
x"8EF171BA",
x"90AE7220",
x"92747262",
x"942A727C",
x"95B97274",
x"97147251",
x"98327223",
x"991271FB",
x"99B871E8",
x"9A2971F9",
x"9A6B7236",
x"9A87729D",
x"9A7D7327",
x"9A4F73C8",
x"99FE746E",
x"998E7502",
x"99037576",
x"986375BE",
x"97BF75D5",
x"972775C1",
x"96AC7590",
x"96637552",
x"965C751F",
x"969F7506",
x"972E751A",
x"98017560",
x"990875D5",
x"9A317671",
x"9B5D7725",
x"9C7877DB",
x"9D6C7883",
x"9E29790E",
x"9EA7796E",
x"9EE379A0",
x"9EE279A6",
x"9EA77986",
x"9E367946",
x"9D9578ED",
x"9CC3787E",
x"9BB977F9",
x"9A74775A",
x"98EE769C",
x"972475B7",
x"951774A7",
x"92D5736C",
x"906E7209",
x"8E00708C",
x"8BA46F02",
x"897E6D82",
x"87AA6C1E",
x"86416AEF",
x"85506A04",
x"84DF6968",
x"84E76921",
x"855B692B",
x"86206980",
x"871B6A11",
x"88326ACF",
x"89486BA8",
x"8A436C8C",
x"8B146D69",
x"8BAF6E35",
x"8C146EE5",
x"8C436F72",
x"8C436FD8",
x"8C217014",
x"8BE37027",
x"8B90700F",
x"8B276FCB",
x"8AA56F5B",
x"8A006EBF",
x"89256DF5",
x"88036CFC",
x"86866BD5",
x"849A6A7F",
x"823768FF",
x"7F596759",
x"7C0B6597",
x"786563C2",
x"748361E8",
x"70916017",
x"6CBD5E5F",
x"69375CD0",
x"662A5B77",
x"63B85A5F",
x"61FC598A",
x"60FB58FD",
x"60B058B2",
x"610958A5",
x"61EB58CD",
x"63315922",
x"64BA599B",
x"66635A32",
x"68175AE4",
x"69C45BB1",
x"6B655C97",
x"6D005D98",
x"6E9D5EB3",
x"704E5FE4",
x"721C6127",
x"7410626D",
x"762E63AF",
x"787064DE",
x"7AC965EC",
x"7D2866D1",
x"7F7C6789",
x"81B26813",
x"83BC6877",
x"859768C4",
x"87426906",
x"88C5694F",
x"8A2C69B2",
x"8B896A3B",
x"8CE66AF5",
x"8E4F6BDF",
x"8FC86CF8",
x"914B6E35",
x"92CC6F8A",
x"943E70E2",
x"958A722A",
x"969F734E",
x"976D743D",
x"97E974E8",
x"9813754B",
x"97F17565",
x"979A753D",
x"972174E7",
x"96AB7475",
x"96577408",
x"964973BB",
x"969D73AA",
x"976773EE",
x"98B57493",
x"9A80759F",
x"9CB87705",
x"9F3F78B4",
x"A1EE7A8B",
x"A4957C65",
x"A7057E1B",
x"A90F7F85",
x"AA948088",
x"AB7D8112",
x"ABC6811B",
x"AB7A80AC",
x"AAB57FD7",
x"A99C7EBC",
x"A85A7D7A",
x"A71B7C33",
x"A6007B05",
x"A5277A0B",
x"A4997950",
x"A45D78DB",
x"A46678AA",
x"A4A478B6",
x"A50478EE",
x"A5717947",
x"A5DE79B4",
x"A6427A29",
x"A6997AA0",
x"A6E77B13",
x"A7327B7F",
x"A7837BE4",
x"A7DD7C40",
x"A8467C91",
x"A8BF7CD6",
x"A9427D0E",
x"A9CC7D39",
x"AA537D56",
x"AAD07D67",
x"AB3B7D6E",
x"AB877D6B",
x"ABAC7D61",
x"ABA17D51",
x"AB597D39",
x"AACC7D14",
x"A9F37CE0",
x"A8CA7C98",
x"A7577C37",
x"A5A37BBF",
x"A3C77B2F",
x"A1DF7A8E",
x"A00F79E7",
x"9E7E7946",
x"9D4F78B7",
x"9C9C784A",
x"9C747803",
x"9CD277E7",
x"9DA277EF",
x"9EC07813",
x"9FFA7841",
x"A11B7868",
x"A1EB7872",
x"A240784E",
x"A1FD77F4",
x"A114775B",
x"9F8D7689",
x"9D7E7583",
x"9B0B7458",
x"985C7317",
x"959571CD",
x"92D87085",
x"90316F45",
x"8DA76E0F",
x"8B2E6CDC",
x"88B26BA6",
x"86206A63",
x"83626910",
x"806C67A7",
x"7D46662D",
x"7A0264AB",
x"76C46334",
x"73BD61DA",
x"712160B8",
x"6F275FE2",
x"6DFC5F6D",
x"6DC15F67",
x"6E825FD8",
x"703A60BB",
x"72D16206",
x"761E63A8",
x"79F0658D",
x"7E11679A",
x"824C69BB",
x"86746BD9",
x"8A666DE6",
x"8E0D6FD9",
x"915A71AF",
x"94507362",
x"96F774FB",
x"99577678",
x"9B8377E1",
x"9D877934",
x"9F707A72",
x"A1487B99",
x"A3157CA5",
x"A4DC7D92",
x"A69C7E5E",
x"A8547F08",
x"AA017F95",
x"AB9C8005",
x"AD1F805E",
x"AE8180A5",
x"AFB680D9",
x"B0B38100",
x"B16E8114",
x"B1DC8114",
x"B1F280FB",
x"B1AF80C3",
x"B10F806A",
x"B0197FF0",
x"AED67F57",
x"AD547EA9",
x"ABAC7DEE",
x"A9EE7D33",
x"A8387C82",
x"A6A17BE8",
x"A53D7B6A",
x"A4217B0B",
x"A3537AC7",
x"A2DA7A99",
x"A2AF7A78",
x"A2C97A5A",
x"A3157A39",
x"A3827A0C",
x"A3FA79D6",
x"A4697998",
x"A4BD7958",
x"A4EC7922",
x"A4EE78FB",
x"A4C378ED",
x"A47078FC",
x"A3FB792A",
x"A36D7974",
x"A2D279D0",
x"A22E7A33",
x"A18A7A96",
x"A0E97AEB",
x"A04D7B2A",
x"9FB97B50",
x"9F2E7B5B",
x"9EB17B51",
x"9E467B36",
x"9DF77B15",
x"9DCF7AF9",
x"9DD77AEB",
x"9E187AF5",
x"9E997B1C",
x"9F5A7B60",
x"A0537BC0",
x"A17A7C34",
x"A2B87CB7",
x"A3F87D3D",
x"A51F7DBA",
x"A6177E25",
x"A6CA7E74",
x"A7327EA5",
x"A7497EB3",
x"A7177EA2",
x"A6AC7E77",
x"A6197E37",
x"A5767DED",
x"A4D27D9F",
x"A4387D51",
x"A3AF7D06",
x"A3327CBF",
x"A2B57C74",
x"A22C7C1E",
x"A18A7BB4",
x"A0C67B32",
x"9FDF7A93",
x"9EE279DE",
x"9DE2791B",
x"9CFD785B",
x"9C5677B3",
x"9C0A773A",
x"9C2F7706",
x"9CD07726",
x"9DE3779D",
x"9F4F7867",
x"A0EB7971",
x"A2847A9F",
x"A3E37BCE",
x"A4D67CDE",
x"A5397DAC",
x"A4FA7E20",
x"A41A7E30",
x"A2AE7DDE",
x"A0DC7D33",
x"9ECF7C47",
x"9CB27B2F",
x"9AA67A03",
x"98BC78D4",
x"96EE77A6",
x"95277674",
x"933C7531",
x"90FE73CB",
x"8E3B7229",
x"8ACF703B",
x"86A86DF9",
x"81CF6B65",
x"7C686891",
x"76B0659A",
x"70F762A5",
x"6B985FDF",
x"66EE5D6D",
x"63405B74",
x"60C85A0B",
x"5FA1593F",
x"5FC8590B",
x"611F5964",
x"636D5A2F",
x"666F5B53",
x"69D85CAF",
x"6D5F5E28",
x"70C45FA7",
x"73D2611A",
x"766F6277",
x"788963B7",
x"7A2364D8",
x"7B4C65DB",
x"7C1966BF",
x"7CA36786",
x"7D036830",
x"7D5068BB",
x"7D9B692A",
x"7DF0697C",
x"7E5569B5",
x"7ECF69DC",
x"7F5969F6",
x"7FF36A0D",
x"80966A2A",
x"81396A54",
x"81D56A8D",
x"82606AD8",
x"82D36B31",
x"83246B92",
x"834C6BEC",
x"83486C38",
x"83156C68",
x"82B56C70",
x"822B6C4E",
x"81806BFD",
x"80BE6B82",
x"7FEF6AE3",
x"7F216A30",
x"7E5F6975",
x"7DB468BF",
x"7D286820",
x"7CC4679E",
x"7C876741",
x"7C766709",
x"7C8E66F0",
x"7CC966EF",
x"7D2366FA",
x"7D936707",
x"7E14670E",
x"7E9E6707",
x"7F2A66F5",
x"7FB466D9",
x"803866BC",
x"80B166AB",
x"811E66B0",
x"817A66D1",
x"81C36716",
x"81F7677C",
x"82116800",
x"82136894",
x"81F9692B",
x"81CB69B5",
x"818D6A26",
x"814B6A72",
x"81146A99",
x"80F76A9D",
x"81066A8A",
x"814E6A6D",
x"81D86A5C",
x"82AA6A63",
x"83BE6A94",
x"85096AF6",
x"86776B89",
x"87F46C48",
x"89646D28",
x"8AB16E16",
x"8BC66F00",
x"8C986FD5",
x"8D217083",
x"8D627102",
x"8D65714B",
x"8D35715F",
x"8CE07144",
x"8C747100",
x"8BFA70A3",
x"8B767035",
x"8AE96FC3",
x"8A526F54",
x"89AF6EEE",
x"88FE6E94",
x"88416E4A",
x"87796E0C",
x"86B46DD9",
x"85FA6DB0",
x"855D6D8A",
x"84E76D6C",
x"84A76D52",
x"84A06D41",
x"84D06D37",
x"85326D38",
x"85B86D44",
x"864E6D59",
x"86DC6D78",
x"874D6D97",
x"87916DB1",
x"879A6DC1",
x"87626DBD",
x"86ED6D9E",
x"86486D66",
x"85866D14",
x"84BC6CAE",
x"84016C38",
x"83666BBE",
x"82F06B45",
x"829E6AD2",
x"825F6A63",
x"821369EF",
x"81906966",
x"80AA68B5",
x"7F3067C5",
x"7CFA667F",
x"79F064D3",
x"761062B9",
x"71696038",
x"6C285D64",
x"668F5A5D",
x"60EC5750",
x"5B9C5471",
x"56F351F1",
x"53405002",
x"50BA4EC3",
x"4F804E49",
x"4F994E95",
x"50E94F93",
x"53435126",
x"5665531C",
x"5A055547",
x"5DD75775",
x"6197597A",
x"65105B36",
x"68195C9A",
x"6A9C5D9F",
x"6C935E52",
x"6E075EC2",
x"6F0C5F08",
x"6FB75F3F",
x"70235F7A",
x"70695FC8",
x"709E6031",
x"70D260B4",
x"710E6146",
x"715961DA",
x"71B0625F",
x"721062C5",
x"72726300",
x"72CC6304",
x"731762D0",
x"73496268",
x"735F61D0",
x"73536118",
x"732A604D",
x"72E55F7D",
x"72905EB3",
x"72325DFD",
x"71DB5D5F",
x"718E5CDD",
x"71565C7D",
x"71345C39",
x"71285C12",
x"712E5C04",
x"713E5C0A",
x"71515C22",
x"715E5C4B",
x"71615C80",
x"71565CC3",
x"713F5D11",
x"71215D6C",
x"71005DCF",
x"70E35E39",
x"70CF5EAB",
x"70C75F1F",
x"70CE5F92",
x"70DF6004",
x"70F9606E",
x"711660D0",
x"71316128",
x"71476173",
x"715261B4",
x"715361E8",
x"714B620E",
x"71386229",
x"711D6238",
x"70FD6239",
x"70DB622D",
x"70B86211",
x"709A61E9",
x"708461B2",
x"707D616F",
x"708C611F",
x"70B760CB",
x"71046072",
x"7177601A",
x"72115FC8",
x"72CE5F80",
x"73A55F49",
x"748A5F24",
x"756F5F15",
x"763F5F1E",
x"76EC5F41",
x"77665F7D",
x"77A75FD2",
x"77AA603B",
x"777060B5",
x"7706613B",
x"767561C5",
x"75CC624C",
x"752062C6",
x"7479632F",
x"73E56380",
x"736963B4",
x"730963C9",
x"72C163C4",
x"728E63A5",
x"726C6374",
x"72556339",
x"724462FA",
x"723762BF",
x"722D628B",
x"72266266",
x"7223624C",
x"7227623E",
x"72316237",
x"72456234",
x"72616231",
x"72806228",
x"72A4621B",
x"72C86206",
x"72E661ED",
x"72FD61D3",
x"730961BB",
x"730461AB",
x"72EF61A2",
x"72C761A5",
x"728761AE",
x"723061B8",
x"71BB61BB",
x"712861AD",
x"7070617D",
x"6F8F6124",
x"6E806094",
x"6D3F5FC6",
x"6BC85EB8",
x"6A1A5D6C",
x"68385BEA",
x"66275A40",
x"63F25880",
x"61A956BF",
x"5F5F5514",
x"5D2D5393",
x"5B305253",
x"5982515E",
x"583B50C4",
x"57735085",
x"573750A2",
x"57885111",
x"586451C7",
x"59B752B5",
x"5B6B53C7",
x"5D5F54EE",
x"5F705615",
x"617D572E",
x"6369582E",
x"651E590B",
x"668F59C5",
x"67BA5A5A",
x"68A45AD3",
x"695C5B36",
x"69F35B8E",
x"6A7A5BE3",
x"6B005C40",
x"6B8E5CAC",
x"6C2A5D2C",
x"6CCF5DC3",
x"6D765E70",
x"6E145F2E",
x"6EA05FF7",
x"6F0F60C3",
x"6F586188",
x"6F7C623E",
x"6F7A62D5",
x"6F596345",
x"6F1E6386",
x"6ED26391",
x"6E7A6365",
x"6E1E6301",
x"6DC4626F",
x"6D6E61B7",
x"6D2460E7",
x"6CEB6015",
x"6CC85F50",
x"6CC15EAB",
x"6CDB5E33",
x"6D175DF3",
x"6D735DEC",
x"6DE95E1C",
x"6E6D5E7A",
x"6EF35EF7",
x"6F695F83",
x"6FC5600E",
x"6FFF608B",
x"701060EC",
x"7001612E",
x"6FDE6150",
x"6FB56158",
x"6F9A614B",
x"6F9B6137",
x"6FC56122",
x"70196117",
x"70916118",
x"71206129",
x"71B16148",
x"7231616D",
x"728C6193",
x"72B861B2",
x"72B161C6",
x"727D61CE",
x"722E61C6",
x"71D661B5",
x"718E61A1",
x"716B6190",
x"71776188",
x"71BB6193",
x"723261B1",
x"72D161E3",
x"73836225",
x"74356273",
x"74D462C4",
x"754C630D",
x"75976349",
x"75B16373",
x"759B6387",
x"755C6386",
x"74FF6376",
x"748A635C",
x"74096341",
x"737C632A",
x"72EB631D",
x"7252631D",
x"71B86328",
x"711B633C",
x"70806353",
x"6FEF6365",
x"6F6D636A",
x"6F04635F",
x"6EBF633E",
x"6EA36306",
x"6EB162B9",
x"6EE9625D",
x"6F4761F3",
x"6FBC6183",
x"70416110",
x"70C2609E",
x"7135602F",
x"718C5FC6",
x"71BE5F60",
x"71C75EFD",
x"71A75E9B",
x"71615E3C",
x"70FC5DE2",
x"70805D8D",
x"6FF65D3F",
x"6F665CFD",
x"6ED25CCB",
x"6E3B5CA5",
x"6DA05C90",
x"6CF65C84",
x"6C375C7E",
x"6B5B5C76",
x"6A5C5C60",
x"693A5C39",
x"67FC5BF7",
x"66B35B98",
x"65765B21",
x"64655A97",
x"63A15A0A",
x"634B598B",
x"637F5932",
x"644D5915",
x"65BB5947",
x"67C159D9",
x"6A475ACD",
x"6D2B5C22",
x"70485DC9",
x"73755FAE",
x"768B61B7",
x"797563C5",
x"7C2465C1",
x"7E9D6794",
x"80EC6937",
x"832E6AA8",
x"85806BF2",
x"87FE6D23",
x"8ABF6E52",
x"8DD26F92",
x"913270F2",
x"94D37278",
x"989A7421",
x"9C6775E4",
x"A01577AA",
x"A381795D",
x"A68E7AE5",
x"A9297C2F",
x"AB497D2C",
x"ACF07DDA",
x"AE257E3C",
x"AEFE7E60",
x"AF8B7E56",
x"AFE07E32",
x"B00E7E07",
x"B01F7DE3",
x"B0197DCF",
x"B0007DCF",
x"AFCF7DE0",
x"AF7F7DFC",
x"AF0F7E1C",
x"AE787E35",
x"ADB97E40",
x"ACD47E37",
x"ABCC7E16",
x"AAA87DE0",
x"A9757D95",
x"A83F7D3C",
x"A7147CD9",
x"A6047C75",
x"A5217C18",
x"A47B7BCC",
x"A4227B99",
x"A4227B85",
x"A4857B99",
x"A54C7BD7",
x"A6707C3F",
x"A7E37CD0",
x"A98E7D7F",
x"AB537E44",
x"AD0B7F0C",
x"AE947FCA",
x"AFCF806B",
x"B09F80DE",
x"B0F88118",
x"B0DE8114",
x"B06080D3",
x"AF9B805D",
x"AEB67FC3",
x"ADE07F1F",
x"AD407E88",
x"ACFE7E15",
x"AD297DDE",
x"ADCD7DF2",
x"AEDC7E53",
x"B03C7EFA",
x"B1C67FD4",
x"B34C80CC",
x"B49F81BD",
x"B5988288",
x"B616830E",
x"B6098338",
x"B56E82FD",
x"B452825C",
x"B2CC8163",
x"B0FD802C",
x"AF087ED7",
x"AD127D82",
x"AB3B7C4E",
x"A9947B53",
x"A8297A9D",
x"A6FD7A32",
x"A6077A05",
x"A5357A08",
x"A4747A20",
x"A3B27A36",
x"A2DD7A33",
x"A1EB7A05",
x"A0DA79A5",
x"9FB17913",
x"9E7B785B",
x"9D4F778B",
x"9C3F76B9",
x"9B5F75F9",
x"9ABC7562",
x"9A6074FE",
x"9A4974D2",
x"9A6D74E2",
x"9AB87520",
x"9B15757F",
x"9B6A75EA",
x"9BA1764E",
x"9BA57697",
x"9B6E76B7",
x"9AF776A3",
x"9A467657",
x"996475D8",
x"9862752D",
x"97487461",
x"9622737E",
x"94EF728F",
x"93A57199",
x"9235709D",
x"90866F94",
x"8E796E78",
x"8BF46D3A",
x"88E36BCE",
x"853A6A2B",
x"8101684E",
x"7C4F663B",
x"775163FF",
x"723B61B1",
x"6D555F6D",
x"68E35D56",
x"65275B8A",
x"62565A26",
x"6096593C",
x"5FF358D4",
x"606458EB",
x"61C8596E",
x"63F25A45",
x"66A45B4F",
x"69A05C6D",
x"6CAA5D83",
x"6F915E7A",
x"72355F49",
x"74825FF3",
x"76756081",
x"781D6108",
x"798E619F",
x"7AE5625A",
x"7C38634C",
x"7D9E647C",
x"7F2465E6",
x"80CF6780",
x"82976934",
x"84716AE5",
x"86486C78",
x"88066DCF",
x"89956EDB",
x"8AE06F8A",
x"8BD86FDF",
x"8C706FDC",
x"8CA86F92",
x"8C816F14",
x"8C096E79",
x"8B4E6DD5",
x"8A666D3D",
x"896C6CBD",
x"88796C5C",
x"87A76C21",
x"87066C06",
x"86A76C04",
x"868A6C13",
x"86AB6C27",
x"86F96C35",
x"875C6C38",
x"87BC6C2A",
x"87FD6C07",
x"88086BD4",
x"87D36B96",
x"87596B55",
x"86A46B1D",
x"85CC6AF9",
x"84ED6AF2",
x"842B6B0D",
x"83A46B4E",
x"83726BB1",
x"839F6C2E",
x"842F6CBA",
x"85116D47",
x"862A6DC5",
x"87596E2A",
x"88766E6B",
x"89626E83",
x"89FE6E73",
x"8A3F6E3F",
x"8A1E6DF2",
x"89A56D94",
x"88E96D30",
x"88016CCF",
x"870A6C75",
x"861A6C26",
x"85446BDE",
x"84916B9C",
x"84066B57",
x"839A6B0C",
x"83456AB5",
x"82F76A52",
x"82A569E3",
x"8245696C",
x"81D368F5",
x"81526886",
x"80C9682A",
x"804567E9",
x"7FD367C9",
x"7F8067CF",
x"7F5667F9",
x"7F596842",
x"7F8768A4",
x"7FD56910",
x"8035697C",
x"809469DB",
x"80DD6A1E",
x"80FE6A42",
x"80E66A3E",
x"808D6A10",
x"7FF269BC",
x"7F186948",
x"7E1068B5",
x"7CE66810",
x"7BAF675C",
x"7A8266A1",
x"796965E2",
x"78756525",
x"77AA646C",
x"770A63BC",
x"76936318",
x"763C6284",
x"75FD6206",
x"75CE619F",
x"75A56153",
x"75836124",
x"7565610E",
x"754E610D",
x"7547611A",
x"7551612E",
x"7573613E",
x"75AF6145",
x"75FF613B",
x"7658611E",
x"76AB60EA",
x"76E560A2",
x"76EB6046",
x"76A55FDA",
x"76015F60",
x"74F05ED9",
x"736F5E45",
x"71825DA5",
x"6F3C5CFD",
x"6CBA5C4D",
x"6A205B9F",
x"67965AFD",
x"65475A6E",
x"63585A05",
x"61E659CC",
x"610959CD",
x"60C45A10",
x"61115A92",
x"61E35B50",
x"631E5C3C",
x"64A35D42",
x"664F5E4D",
x"68005F45",
x"699C6015",
x"6B0D60AE",
x"6C476104",
x"6D426117",
x"6E0760EC",
x"6E9A608E",
x"6F096013",
x"6F5F5F8D",
x"6FA85F0E",
x"6FED5EAB",
x"70315E6E",
x"70725E5C",
x"70AD5E76",
x"70DE5EB2",
x"70FD5F08",
x"710A5F6C",
x"71035FD0",
x"70ED602D",
x"70D2607A",
x"70BB60BB",
x"70B860F0",
x"70D56125",
x"711A6160",
x"718C61AB",
x"7228620D",
x"72E56286",
x"73B56313",
x"748663AB",
x"75456441",
x"75E364C6",
x"7654652D",
x"76966568",
x"76AB6572",
x"76A0654C",
x"768664FF",
x"766F6495",
x"76706425",
x"769763BF",
x"76EF6377",
x"777C635D",
x"783A6377",
x"791D63C9",
x"7A17644E",
x"7B1A64F9",
x"7C1365BB",
x"7CF46683",
x"7DB76741",
x"7E5267E6",
x"7EC56869",
x"7F1168C5",
x"7F3A68FC",
x"7F446911",
x"7F31690C",
x"7F0968F3",
x"7ECC68D1",
x"7E7F68AA",
x"7E276883",
x"7DC8685E",
x"7D696838",
x"7D136814",
x"7CCC67ED",
x"7C9B67C1",
x"7C83678C",
x"7C87674F",
x"7CA5670A",
x"7CD866BC",
x"7D156669",
x"7D566611",
x"7D9065BA",
x"7DB86560",
x"7DC9650A",
x"7DBF64B5",
x"7D9B6465",
x"7D5F6414",
x"7D1063C6",
x"7CB26379",
x"7C4E632D",
x"7BE862E2",
x"7B806298",
x"7B1B6252",
x"7AB76211",
x"7A5161D6",
x"79E861A4",
x"79766179",
x"78FA6153",
x"78756132",
x"77E56113",
x"774F60F2",
x"76B760CB",
x"7623609E",
x"7597606A",
x"751B6032",
x"74B15FF9",
x"745B5FC2",
x"74165F90",
x"73DC5F69",
x"73A75F4C",
x"736F5F3C",
x"732A5F35",
x"72D25F35",
x"72635F38",
x"71DC5F3C",
x"71425F41",
x"709B5F45",
x"6FF05F4C",
x"6F4A5F58",
x"6EAD5F6D",
x"6E1E5F90",
x"6D9D5FBE",
x"6D245FF7",
x"6CAB6035",
x"6C286072",
x"6B94609E",
x"6AE960B2",
x"6A2460A4",
x"694E606A",
x"68736003",
x"67A55F70",
x"66FC5EBB",
x"66905DF3",
x"66795D2B",
x"66CE5C78",
x"679E5BF6",
x"68F65BB9",
x"6AD75BD7",
x"6D3F5C5F",
x"70245D56",
x"73785EBF",
x"7724608E",
x"7B1062B4",
x"7F1E6517",
x"8332679B",
x"872A6A23",
x"8AE96C8D",
x"8E506EC3",
x"914B70AE",
x"93C87247",
x"95BC7386",
x"97297472",
x"98187515",
x"9898757C",
x"98BC75B7",
x"989F75D4",
x"985875DC",
x"97FB75DA",
x"979A75CB",
x"973F75B1",
x"96EE7586",
x"96A97546",
x"966C74EB",
x"96317475",
x"95F773EA",
x"95BE734D",
x"958B72AB",
x"95667212",
x"9556718A",
x"95677124",
x"959C70E5",
x"95F870D1",
x"967670E4",
x"97047116",
x"9790715B",
x"980171A1",
x"983E71DA",
x"982F71F4",
x"97C571E4",
x"96F671A4",
x"95C67137",
x"944570A3",
x"92876FF5",
x"90AB6F3E",
x"8ECB6E8F",
x"8D066DF6",
x"8B6F6D7D",
x"8A146D2D",
x"88FA6D00",
x"881D6CF0",
x"87726CF2",
x"86ED6CF8",
x"86836CF3",
x"862C6CD8",
x"85E66CA0",
x"85AF6C4D",
x"85906BE1",
x"858E6B68",
x"85B16AF2",
x"85FC6A8F",
x"866A6A4F",
x"86F66A3E",
x"87906A65",
x"88256AC4",
x"88A56B57",
x"88FE6C12",
x"89246CE2",
x"89116DB5",
x"88C86E75",
x"884D6F0D",
x"87B16F70",
x"87006F93",
x"864C6F75",
x"85A46F1A",
x"85106E92",
x"84976DEE",
x"843B6D41",
x"83FC6CA3",
x"83D66C23",
x"83C86BCF",
x"83CF6BAD",
x"83EC6BBA",
x"84216BEC",
x"84706C38",
x"84DC6C8D",
x"85636CDB",
x"86066D14",
x"86B96D31",
x"87746D2D",
x"882A6D09",
x"88C66CCB",
x"893E6C7A",
x"89806C23",
x"89886BCC",
x"89536B7D",
x"88E76B3B",
x"88506B0A",
x"879E6AE9",
x"86E36AD8",
x"86326AD2",
x"85986AD5",
x"851E6ADE",
x"84C66AE5",
x"848E6AE8",
x"846D6AE1",
x"84586ACC",
x"84446AA8",
x"84286A75",
x"83FD6A34",
x"83BF69E9",
x"836A6999",
x"82FC6945",
x"826968F2",
x"81A5689A",
x"809B6834",
x"7F3267B4",
x"7D4E6703",
x"7AD1660D",
x"77A764BB",
x"73C962FD",
x"6F4160CC",
x"6A275E2B",
x"64AD5B2E",
x"5F1057F4",
x"599A54AC",
x"54995189",
x"50514EC4",
x"4CFF4C8C",
x"4AC84B08",
x"49BD4A4E",
x"49D44A62",
x"4AEF4B34",
x"4CDF4CA3",
x"4F6B4E85",
x"525250A5",
x"555C52D0",
x"585754DC",
x"5B1956A6",
x"5D8A581E",
x"5FA4593C",
x"61655A0A",
x"62DB5A97",
x"64135AF8",
x"65235B46",
x"661A5B92",
x"67065BE9",
x"67EF5C4F",
x"68D65CC3",
x"69BA5D3C",
x"6A915DAE",
x"6B535E0B",
x"6BF95E48",
x"6C7A5E5D",
x"6CD55E49",
x"6D0C5E10",
x"6D275DBD",
x"6D315D62",
x"6D375D0D",
x"6D495CD2",
x"6D725CBD",
x"6DB85CDD",
x"6E1B5D31",
x"6E965DB1",
x"6F1B5E53",
x"6F9B5F03",
x"70015FA8",
x"703B602E",
x"703A6080",
x"6FF3608E",
x"6F656058",
x"6E965FDD",
x"6D905F2C",
x"6C665E5A",
x"6B2D5D7E",
x"69F95CB2",
x"68DF5C0A",
x"67EE5B94",
x"67315B59",
x"66AB5B56",
x"665E5B80",
x"663F5BC8",
x"664A5C1A",
x"666C5C60",
x"669B5C8E",
x"66CC5C98",
x"66F55C7B",
x"670F5C3D",
x"67195BEA",
x"67165B91",
x"670A5B45",
x"67005B14",
x"66FF5B0B",
x"67105B33",
x"673B5B8B",
x"67855C0B",
x"67EE5CA8",
x"68755D52",
x"69145DF8",
x"69C85E8E",
x"6A8C5F0A",
x"6B595F64",
x"6C2B5FA2",
x"6D025FC6",
x"6DD65FD9",
x"6EAA5FE6",
x"6F765FF3",
x"70376007",
x"70E36022",
x"71756042",
x"71E1605F",
x"721E6072",
x"722B6073",
x"7209605D",
x"71BC6032",
x"71515FF4",
x"70D65FAF",
x"705F5F6E",
x"6FFD5F43",
x"6FBE5F38",
x"6FAD5F56",
x"6FCB5FA2",
x"7014601A",
x"707F60AF",
x"70FC6156",
x"717D61F9",
x"71F06284",
x"724B62E9",
x"72846317",
x"72966307",
x"728262BB",
x"724B6238",
x"71F56187",
x"718760B8",
x"71065FDA",
x"70775EFC",
x"6FDF5E2B",
x"6F445D6E",
x"6EA85CCD",
x"6E145C48",
x"6D8F5BDD",
x"6D1E5B88",
x"6CC75B46",
x"6C8A5B11",
x"6C665AE3",
x"6C515AB9",
x"6C385A90",
x"6C0A5A63",
x"6BB05A30",
x"6B0E59F4",
x"6A1659A9",
x"68B5594A",
x"66EC58D3",
x"64C25840",
x"624B578F",
x"5FA456C0",
x"5CF555D9",
x"5A6654DE",
x"582153E1",
x"564E52EE",
x"55065218",
x"545E5171",
x"545C510B",
x"54FF50F1",
x"5637512F",
x"57EC51C3",
x"5A0552AB",
x"5C6253D9",
x"5EE2553C",
x"616956BF",
x"63DC584C",
x"662759CA",
x"68385B2B",
x"6A0A5C5F",
x"6B9A5D60",
x"6CEE5E2F",
x"6E0D5ED3",
x"6F075F58",
x"6FEC5FC9",
x"70C86037",
x"71A660AB",
x"728C612B",
x"737C61B9",
x"74726252",
x"756562EC",
x"764A637C",
x"771963FA",
x"77C86460",
x"785664AA",
x"78C564D9",
x"791A64F7",
x"7960650B",
x"79A46521",
x"79EC6541",
x"7A3F6570",
x"7A9D65AD",
x"7AFD65F0",
x"7B566632",
x"7B986666",
x"7BB7667F",
x"7BA46676",
x"7B5C6646",
x"7AE065F6",
x"7A3D6591",
x"79806528",
x"78C164CC",
x"781A6491",
x"77A06487",
x"776664B5",
x"777A651D",
x"77E265B8",
x"789A6679",
x"79986751",
x"7ACF682D",
x"7C2B68FD",
x"7D9569B4",
x"7EF96A4C",
x"80446AC5",
x"81636B21",
x"824F6B68",
x"82FE6BA0",
x"83726BD4",
x"83AE6C07",
x"83BC6C3F",
x"83AD6C7C",
x"838E6CBA",
x"83736CFA",
x"836D6D38",
x"83876D72",
x"83CC6DA9",
x"843F6DDC",
x"84E06E10",
x"85A46E43",
x"86836E76",
x"876C6EA9",
x"88506ED7",
x"89216EFA",
x"89D06F0F",
x"8A566F0C",
x"8AAA6EEE",
x"8AC96EB3",
x"8AB56E5C",
x"8A706DF0",
x"8A016D76",
x"896C6CF5",
x"88B76C75",
x"87EA6BF9",
x"87086B87",
x"861A6B1A",
x"85216AB0",
x"84206A41",
x"831E69C7",
x"82206941",
x"812E68AE",
x"80516814",
x"7F946780",
x"7F0466FD",
x"7EAB669A",
x"7E936663",
x"7EBC665C",
x"7F286687",
x"7FC866D8",
x"808C673E",
x"815B67A4",
x"821867F0",
x"82AA6810",
x"82F467F2",
x"82E66791",
x"827366F3",
x"81A06624",
x"8074653B",
x"7F04644F",
x"7D666377",
x"7BB162C6",
x"79F46241",
x"783A61E8",
x"767F61A9",
x"74BA6176",
x"72DC6131",
x"70D160C3",
x"6E8C601E",
x"6C075F39",
x"694C5E1B",
x"66765CD3",
x"63AE5B81",
x"61275A45",
x"5F1D5945",
x"5DC8589F",
x"5D585870",
x"5DEC58C3",
x"5F8D5997",
x"62305AE3",
x"65B35C90",
x"69E35E83",
x"6E8360A2",
x"735362D0",
x"781A64FC",
x"7CA16713",
x"80C8690D",
x"84766AEB",
x"87A56CAA",
x"8A596E4B",
x"8C9A6FCD",
x"8E7A712D",
x"90067268",
x"914F7375",
x"92607450",
x"934674F6",
x"940B756B",
x"94B875B4",
x"955675DE",
x"95F075F9",
x"968D7615",
x"97357641",
x"97ED768B",
x"98B276F5",
x"9981777F",
x"9A527820",
x"9B1A78CE",
x"9BCF797B",
x"9C647A16",
x"9CD67A96",
x"9D1E7AF5",
x"9D3D7B2F",
x"9D397B46",
x"9D1A7B3E",
x"9CE77B20",
x"9CAC7AEF",
x"9C707AAF",
x"9C397A61",
x"9C087A03",
x"9BDD7995",
x"9BB67910",
x"9B8D7878",
x"9B5C77CA",
x"9B1A770D",
x"9AC07647",
x"9A4D7582",
x"99BE74C7",
x"990E741F",
x"98457390",
x"9767731F",
x"967D72CA",
x"9590728D",
x"94AA7264",
x"93D27244",
x"93117229",
x"92677209",
x"91D371E1",
x"914F71AF",
x"90D27174",
x"90557130",
x"8FCC70E6",
x"8F34709D",
x"8E887057",
x"8DCD7017",
x"8D0D6FDF",
x"8C4E6FB4",
x"8B9F6F97",
x"8B106F8A",
x"8AA56F92",
x"8A696FAE",
x"8A596FE1",
x"8A737027",
x"8AAC7082",
x"8AFA70EB",
x"8B50715E",
x"8BA471D1",
x"8BEC723A",
x"8C257293",
x"8C5272D2",
x"8C7172F1",
x"8C8E72EF",
x"8CAC72CD",
x"8CD37290",
x"8D087243",
x"8D4F71EE",
x"8DA7719C",
x"8E0D7157",
x"8E7D7127",
x"8EF0710F",
x"8F5D710C",
x"8FBE7119",
x"9008712D",
x"9039713E",
x"90487143",
x"90327133",
x"8FF7710C",
x"8F9770CD",
x"8F127079",
x"8E70701D",
x"8DB56FBE",
x"8CE76F68",
x"8C116F24",
x"8B386EF6",
x"8A696EDF",
x"89AE6EDC",
x"89116EE9",
x"889E6F02",
x"88636F1E",
x"88676F40",
x"88B26F65",
x"89426F92",
x"8A136FCA",
x"8B0E7010",
x"8C1A7064",
x"8D0D70BD",
x"8DB97108",
x"8DEA7131",
x"8D6D7119",
x"8C18709F",
x"89CF6FA9",
x"868B6E21",
x"825D6C02",
x"7D6F6955",
x"77FF6635",
x"725C62D2",
x"6CE25F63",
x"67E65C28",
x"63B8595F",
x"6096573A",
x"5EA355E4",
x"5DEC556B",
x"5E6355CD",
x"5FE656F1",
x"624258AE",
x"653E5AD2",
x"689B5D25",
x"6C265F73",
x"6FAD6191",
x"730C635F",
x"762864CC",
x"78EF65D5",
x"7B556681",
x"7D5566E2",
x"7EEC670B",
x"80186713",
x"80E0670A",
x"814B6700",
x"816666FF",
x"8145670B",
x"80FD6727",
x"80AA6752",
x"80656789",
x"804567C9",
x"805C6813",
x"80B16865",
x"814268BB",
x"82036917",
x"82E26976",
x"83C569D4",
x"84946A2B",
x"85366A7A",
x"859B6ABA",
x"85B56AE5",
x"85846AF9",
x"850B6AF3",
x"84566AD5",
x"83766A9E",
x"827C6A55",
x"817A69FD",
x"8084699D",
x"7FAA6938",
x"7EF768D8",
x"7E776881",
x"7E30683B",
x"7E25680A",
x"7E5667F5",
x"7EBF67FF",
x"7F56682A",
x"8011687A",
x"80DD68EB",
x"81AE6976",
x"826F6A16",
x"83136ABF",
x"83906B65",
x"83DF6BFA",
x"84046C73",
x"84066CC8",
x"83F26CF2",
x"83D86CF2",
x"83C96CCD",
x"83D56C8A",
x"840A6C3B",
x"846F6BEC",
x"85046BAD",
x"85CC6B8F",
x"86BC6B99",
x"87CC6BD2",
x"88EF6C3A",
x"8A176CCD",
x"8B356D7C",
x"8C3B6E38",
x"8D1D6EF2",
x"8DCF6F94",
x"8E457010",
x"8E7A7055",
x"8E6A705F",
x"8E15702A",
x"8D806FBE",
x"8CB56F27",
x"8BC46E78",
x"8AB96DC2",
x"89A86D1E",
x"88A46CA0",
x"87B76C54",
x"86ED6C41",
x"864B6C6C",
x"85CE6CCB",
x"85716D4F",
x"852E6DE6",
x"84F96E79",
x"84C86EF2",
x"84936F3D",
x"84566F4D",
x"84116F17",
x"83C86EA0",
x"837D6DEB",
x"833B6D0A",
x"83046C0F",
x"82E06B0F",
x"82CE6A20",
x"82CC6956",
x"82D368C1",
x"82DE686B",
x"82DF6854",
x"82CF6879",
x"82A768D1",
x"825F694B",
x"81F769D5",
x"81746A5B",
x"80DC6ACB",
x"80376B16",
x"7F906B30",
x"7EEF6B11",
x"7E596ABB",
x"7DD06A32",
x"7D53697C",
x"7CD968A4",
x"7C5667B4",
x"7BBE66BA",
x"7B0265BE",
x"7A1A64CC",
x"78FF63E9",
x"77B1631F",
x"763A6273",
x"74AB61EA",
x"731D618A",
x"71B06158",
x"70876156",
x"6FCA618B",
x"6F9B61F6",
x"70196298",
x"71526370",
x"734F647C",
x"760465B5",
x"79586719",
x"7D23689D",
x"81316A3D",
x"854B6BEB",
x"89386DA0",
x"8CC66F51",
x"8FCF70F2",
x"923F7276",
x"941173D4",
x"95557502",
x"962775FB",
x"96AF76B9",
x"9715773E",
x"97817790",
x"980E77B6",
x"98C877B9",
x"99AF77A3",
x"9AB27781",
x"9BB8775A",
x"9CA27734",
x"9D537715",
x"9DB376FC",
x"9DB976EB",
x"9D6476E0",
x"9CC376DB",
x"9BED76DB",
x"9AFE76E1",
x"9A1276EC",
x"994376FF",
x"989B7715",
x"9821772C",
x"97CD773E",
x"97947747",
x"9760773D",
x"9725771D",
x"96D376E5",
x"96667697",
x"95DF763C",
x"954B75DC",
x"94B9758C",
x"943C7555",
x"93E37546",
x"93BC7567",
x"93CB75B7",
x"940B7633",
x"947476CD",
x"94F4776F",
x"957B7808",
x"95F67882",
x"965778CB",
x"969A78DA",
x"96BC78AA",
x"96C87840",
x"96C577A2",
x"96C376E1",
x"96D3760F",
x"9700753E",
x"9750747F",
x"97C973E2",
x"98697374",
x"9925733D",
x"99F47343",
x"9AC67389",
x"9B8E740C",
x"9C3B74C3",
x"9CBF75A3",
x"9D10769C",
x"9D287798",
x"9D04787F",
x"9CA4793E",
x"9C1079C3",
x"9B4C79FC",
x"9A6979E5",
x"996F7982",
x"986C78DD",
x"976C7803",
x"9673770D",
x"958A7610",
x"94AF751C",
x"93E1743E",
x"931A737E",
x"925572D8",
x"918A724A",
x"90B571C8",
x"8FD5714B",
x"8EEA70CB",
x"8DFC7045",
x"8D116FBD",
x"8C316F37",
x"8B696EBD",
x"8AC16E57",
x"8A3F6E0F",
x"89EA6DE6",
x"89C26DDC",
x"89C36DE9",
x"89E76E03",
x"8A256E1D",
x"8A6F6E2A",
x"8AB86E20",
x"8AF16DF6",
x"8B106DAD",
x"8B096D47",
x"8AD96CCF",
x"8A7C6C4E",
x"89F76BD2",
x"894E6B68",
x"88886B16",
x"87AE6AE2",
x"86C26AC8",
x"85C56AC4",
x"84AF6AC7",
x"83776ABF",
x"820A6A9A",
x"80556A44",
x"7E4469A8",
x"7BCB68BB",
x"78E26779",
x"759365E2",
x"71ED6403",
x"6E1761F0",
x"6A385FC5",
x"66865D9F",
x"63345BA1",
x"607359E6",
x"5E6B5884",
x"5D33578C",
x"5CD15705",
x"5D3B56EB",
x"5E595732",
x"600757CA",
x"6217589F",
x"645E599C",
x"66B75AAC",
x"69035BC2",
x"6B345CCD",
x"6D3F5DCC",
x"6F2E5EB8",
x"710C5F92",
x"72E56060",
x"74C96127",
x"76C161ED",
x"78CE62B8",
x"7AE8638B",
x"7D03646D",
x"7F0B655F",
x"80EC665B",
x"8294675F",
x"83F26863",
x"84FD695C",
x"85B56A3E",
x"861D6AFF",
x"863F6B94",
x"86286BF9",
x"85E76C2A",
x"858A6C2B",
x"851E6C03",
x"84AB6BBB",
x"84386B62",
x"83CB6B02",
x"83656AA4",
x"83096A4F",
x"82B56A03",
x"826D69BE",
x"822E6979",
x"81FA692D",
x"81D068CF",
x"81B1685F",
x"819B67DB",
x"81906745",
x"819366A8",
x"81A46610",
x"81C8658D",
x"8201652B",
x"825364F9",
x"82BC64FC",
x"8339653A",
x"83C165AB",
x"8449664B",
x"84C6670A",
x"852767DC",
x"856368AE",
x"85706975",
x"854E6A26",
x"85006AB8",
x"84956B2D",
x"841E6B84",
x"83AF6BC5",
x"835D6BF8",
x"833E6C24",
x"835A6C52",
x"83BE6C89",
x"84636CCB",
x"85446D1D",
x"864F6D7A",
x"87736DE2",
x"88986E4E",
x"89A96EBA",
x"8A936F1C",
x"8B406F70",
x"8BA76FAE",
x"8BBE6FD1",
x"8B806FD1",
x"8AF06FAB",
x"8A156F5C",
x"88FC6EE6",
x"87B16E4B",
x"864B6D92",
x"84DD6CC2",
x"837F6BEC",
x"82436B1C",
x"813E6A5F",
x"807969BF",
x"7FFA6947",
x"7FC168F7",
x"7FC568CE",
x"7FFD68C5",
x"805668D4",
x"80C268EC",
x"812F6907",
x"8194691B",
x"81E86927",
x"8228692B",
x"8258692E",
x"82796935",
x"82936948",
x"82AD696C",
x"82C8699E",
x"82E669DB",
x"83046A17",
x"831E6A45",
x"832B6A54",
x"83276A3A",
x"830769EC",
x"82CE696D",
x"827768C2",
x"820A67FA",
x"81886727",
x"80F9665E",
x"805F65AF",
x"7FBA6528",
x"7F0164C9",
x"7E2D648D",
x"7D2D6460",
x"7BEF6431",
x"7A6663E5",
x"7889636A",
x"765662B2",
x"73DC61BB",
x"7131608E",
x"6E795F3F",
x"6BDE5DE9",
x"698D5CAC",
x"67B35BAB",
x"666E5AFA",
x"65D55AAC",
x"65EB5AC3",
x"66A15B38",
x"67DC5BF4",
x"69755CE0",
x"6B3D5DDD",
x"6D065ED0",
x"6EAB5FA1",
x"70136042",
x"713160AE",
x"720460EA",
x"729E6100",
x"73146100",
x"73836100",
x"74066110",
x"74B2613F",
x"759A619B",
x"76C1622B",
x"782462EF",
x"79B763E6",
x"7B686507",
x"7D236648",
x"7ED6679D",
x"807068F6",
x"81E86A42",
x"83386B73",
x"84636C79",
x"856F6D48",
x"86636DDB",
x"874B6E2E",
x"882F6E47",
x"89176E31",
x"8A046DFC",
x"8AF36DBA",
x"8BE06D7F",
x"8CC16D5C",
x"8D8B6D5F",
x"8E356D90",
x"8EB96DEF",
x"8F156E75",
x"8F4B6F16",
x"8F5F6FC4",
x"8F607070",
x"8F58710A",
x"8F56718A",
x"8F6771E6",
x"8F947221",
x"8FE4723B",
x"9059723A",
x"90F07227",
x"91A5720A",
x"927171EB",
x"934B71CD",
x"942671B3",
x"94FA719F",
x"95BC7192",
x"9663718C",
x"96E4718D",
x"973B7196",
x"975F71A7",
x"974F71C1",
x"970D71E5",
x"96A17216",
x"96157255",
x"957A72A3",
x"94E672FF",
x"946D736B",
x"942473E5",
x"9417746E",
x"945274FF",
x"94D27595",
x"95907627",
x"967776B1",
x"97737727",
x"98647783",
x"993277BD",
x"99C677D1",
x"9A1277C1",
x"9A147792",
x"99D2774A",
x"995A76F8",
x"98C676A7",
x"982E7665",
x"97A8763A",
x"97457627",
x"970B762F",
x"96F87647",
x"96FB7661",
x"97017671",
x"96EA7662",
x"969E762A",
x"960775BD",
x"9518751A",
x"93D67443",
x"924C7344",
x"909A722D",
x"8EE07110",
x"8D497002",
x"8C006F14",
x"8B226E58",
x"8AC66DD7",
x"8AF36D94",
x"8B9D6D92",
x"8CAC6DC7",
x"8DFC6E2A",
x"8F636EAD",
x"90B96F43",
x"91D96FD9",
x"92AB7065",
x"932470DB",
x"93437135",
x"931B716E",
x"92BF7186",
x"92467180",
x"91C6715F",
x"91467126",
x"90C270D5",
x"90257069",
x"8F4D6FDB",
x"8E126F1E",
x"8C486E27",
x"89C86CE8",
x"867C6B58",
x"82666972",
x"7DA0673C",
x"785964C8",
x"72DC622F",
x"6D805F98",
x"68A35D29",
x"64975B10",
x"61A45970",
x"5FF85869",
x"5FA1580B",
x"60905859",
x"629C5942",
x"65875AAF",
x"69095C7D",
x"6CD55E81",
x"70AD6095",
x"74566297",
x"77B0646D",
x"7AA56607",
x"7D356760",
x"7F666879",
x"8145695B",
x"82E26A0F",
x"84486AA0",
x"85816B16",
x"86916B76",
x"877C6BC4",
x"88416BFD",
x"88E26C26",
x"89646C3D",
x"89D06C47",
x"8A2E6C4A",
x"8A896C4D",
x"8AE66C55",
x"8B4B6C69",
x"8BB56C8C",
x"8C1E6CB8",
x"8C7D6CEB",
x"8CC36D17",
x"8CE66D34",
x"8CDD6D38",
x"8CA16D1C",
x"8C356CDF",
x"8B9B6C83",
x"8ADF6C13",
x"8A0B6B99",
x"892D6B23",
x"884C6ABB",
x"87746A6C",
x"86AA6A37",
x"85F36A1C",
x"85526A14",
x"84CC6A19",
x"84666A20",
x"84276A23",
x"84176A20",
x"843E6A1A",
x"84A46A17",
x"854E6A23",
x"863C6A48",
x"876C6A91",
x"88D06B09",
x"8A5F6BB1",
x"8C036C87",
x"8DA76D85",
x"8F396E9D",
x"90A86FC3",
x"91E370E6",
x"92E371FE",
x"93A172FE",
x"942273E1",
x"946974A1",
x"9481753E",
x"947675B9",
x"9452760D",
x"9422763E",
x"93F0764A",
x"93C0762F",
x"939575EE",
x"93717589",
x"93527506",
x"932F746E",
x"930A73CD",
x"92DA732F",
x"92A272A4",
x"925F723A",
x"921471F9",
x"91C971E9",
x"91847209",
x"914F7251",
x"913172B7",
x"912E732B",
x"9149739F",
x"91837400",
x"91D07443",
x"922C745F",
x"928A7451",
x"92DD741C",
x"931A73C6",
x"93387355",
x"933172D8",
x"9304725A",
x"92B471E2",
x"92487179",
x"91C97123",
x"913E70E2",
x"90B270B5",
x"902B709C",
x"8FAB708F",
x"8F35708D",
x"8EC57090",
x"8E597097",
x"8DEF70A0",
x"8D8670AA",
x"8D2170B9",
x"8CC970CF",
x"8C9070F6",
x"8C867133",
x"8CBF718D",
x"8D527209",
x"8E4672A9",
x"8FA17368",
x"9152743B",
x"93397510",
x"952975D0",
x"96E3765D",
x"981F7696",
x"98977662",
x"980E75A7",
x"9659745B",
x"936A727B",
x"8F527014",
x"8A426D47",
x"848E6A38",
x"7E9E671A",
x"78E56421",
x"73D3617E",
x"6FCF5F5C",
x"6D1D5DD9",
x"6BE55D06",
x"6C265CDF",
x"6DBB5D59",
x"70635E59",
x"73CB5FBE",
x"77946163",
x"7B69632A",
x"7F0464F3",
x"823766B0",
x"84E76854",
x"871D69DE",
x"88EC6B55",
x"8A796CC4",
x"8BF06E34",
x"8D7B6FB0",
x"8F387140",
x"913B72E5",
x"9387749A",
x"9617765B",
x"98D3781B",
x"9BA279CA",
x"9E647B5E",
x"A0FD7CC6",
x"A3537DF8",
x"A5537EEA",
x"A6F17F98",
x"A82C8001",
x"A9048026",
x"A982800F",
x"A9B27FC6",
x"A99F7F53",
x"A9577EC7",
x"A8E77E2D",
x"A85A7D94",
x"A7B57D04",
x"A7017C86",
x"A6427C1E",
x"A57A7BCC",
x"A4AC7B8E",
x"A3DD7B5E",
x"A3107B39",
x"A2467B16",
x"A1877AF5",
x"A0D47AD1",
x"A0337AAA",
x"9FA87A84",
x"9F2F7A5E",
x"9ECC7A3E",
x"9E7B7A26",
x"9E3B7A19",
x"9E0A7A18",
x"9DE67A20",
x"9DD07A34",
x"9DC87A51",
x"9DCC7A72",
x"9DDF7A96",
x"9DFB7AB7",
x"9E1F7AD0",
x"9E427ADB",
x"9E597AD1",
x"9E5A7AB0",
x"9E3B7A72",
x"9DF47A19",
x"9D8179A6",
x"9CE77925",
x"9C2F789F",
x"9B6A7825",
x"9AAB77C4",
x"9A087789",
x"9994777E",
x"9959779F",
x"995A77E7",
x"99927844",
x"99ED78A0",
x"9A5278E2",
x"9AA278F2",
x"9AC078C0",
x"9A947840",
x"9A0D7778",
x"99277677",
x"97EA7550",
x"966C7425",
x"94C9730F",
x"9322722A",
x"91977185",
x"90467124",
x"8F417105",
x"8E917116",
x"8E387144",
x"8E2A7178",
x"8E5771A0",
x"8EAE71B3",
x"8F1871AB",
x"8F8A7192",
x"8FF67175",
x"90597165",
x"90B57175",
x"911071B1",
x"91717221",
x"91E072C3",
x"92637389",
x"92FA7464",
x"939F7539",
x"944B75F4",
x"94F0767F",
x"958476D0",
x"95FE76E1",
x"965776B9",
x"96917664",
x"96B575F8",
x"96CD758D",
x"96EC753B",
x"971E7517",
x"9769752A",
x"97CF7578",
x"984075F6",
x"98A27690",
x"98D27729",
x"98A27799",
x"97E677C0",
x"967A7779",
x"944676AD",
x"914C7550",
x"8D9C7366",
x"896A7108",
x"84F46E57",
x"808D6B83",
x"7C8968C7",
x"79376655",
x"76D96463",
x"759B6317",
x"758A6286",
x"769962B5",
x"78A2639A",
x"7B6D651A",
x"7EB46713",
x"82316958",
x"85A46BC2",
x"88DC6E2B",
x"8BB67073",
x"8E277286",
x"902F7458",
x"91E275E4",
x"9356772F",
x"94A87840",
x"95F47920",
x"974C79DB",
x"98BE7A79",
x"9A4C7B04",
x"9BF17B7F",
x"9DA77BF1",
x"9F5D7C5B",
x"A1057CC0",
x"A2917D20",
x"A3F47D7E",
x"A5297DD9",
x"A62B7E33",
x"A6FB7E8E",
x"A79C7EE8",
x"A8187F45",
x"A8787FA5",
x"A8CA800A",
x"A91B8075",
x"A97880E8",
x"A9F18164",
x"AA9181EB",
x"AB5E827D",
x"AC608319",
x"AD9483C3",
x"AEFA8478",
x"B08B8538",
x"B23B8603",
x"B3FE86D4",
x"B5CA87AE",
x"B791888B",
x"B94C896A",
x"BAF18A46",
x"BC7D8B1B",
x"BDEB8BE7",
x"BF3A8CA5",
x"C0678D50",
x"C1708DE6",
x"C24E8E60",
x"C2FF8EBC",
x"C37B8EF9",
x"C3BC8F13",
x"C3BC8F07",
x"C3788ED8",
x"C2F18E86",
x"C22A8E13",
x"C12C8D83",
x"C0058CE0",
x"BEC68C31",
x"BD828B80",
x"BC548AD9",
x"BB4E8A48",
x"BA8889D6",
x"BA0C898B",
x"B9E7896C",
x"BA168977",
x"BA9389A9",
x"BB4E89FB",
x"BC308A62",
x"BD238AD2",
x"BE098B43",
x"BED08BAC",
x"BF638C0B",
x"BFBA8C62",
x"BFD68CB4",
x"BFBD8D0A",
x"BF818D6A",
x"BF328DDC",
x"BEE38E5D",
x"BE9E8EE7",
x"BE6B8F6C",
x"BE438FD3",
x"BE1C9004",
x"BDDE8FE2",
x"BD718F53",
x"BCBC8E4B",
x"BBAB8CC6",
x"BA338AD0",
x"B8568887",
x"B6228614",
x"B3B383A9",
x"B12F817E",
x"AEBF7FC3",
x"AC8F7E9F",
x"AAC57E23",
x"A9787E4F",
x"A8B87F0A",
x"A87B802B",
x"A8B0817D",
x"A93382C2",
x"A9D683C0",
x"AA69844C",
x"AABD8447",
x"AAB283AF",
x"AA308291",
x"A933810E",
x"A7C67F54",
x"A6007D99",
x"A4027C06",
x"A1F07ABD",
x"9FE679CE",
x"9DF77937",
x"9C2678E0",
x"9A66789F",
x"989A784A",
x"969877AD",
x"943B76A2",
x"915A750B",
x"8DE072E1",
x"89CC7030",
x"852F6D17",
x"803969C5",
x"7B2B6672",
x"76506358",
x"71FC60AE",
x"6E7C5E9F",
x"6C0D5D4C",
x"6AD95CC3",
x"6AF25D04",
x"6C4C5E01",
x"6ECE5FA1",
x"724761C8",
x"76806455",
x"7B446727",
x"805B6A20",
x"85976D2A",
x"8AD6702B",
x"8FFE7315",
x"94FB75D7",
x"99C07867",
x"9E437ABC",
x"A2777CD0",
x"A64F7EA0",
x"A9BD802C",
x"ACB58178",
x"AF268288",
x"B10B8366",
x"B2618417",
x"B32B84A3",
x"B3748514",
x"B352856D",
x"B2D985B1",
x"B22385DE",
x"B14C85F7",
x"B06B85F4",
x"AF9185D7",
x"AEC7859B",
x"AE12853D",
x"AD6A84BD",
x"ACC5841B",
x"AC0E8354",
x"AB368268",
x"AA30815B",
x"A8F3802D",
x"A77F7EE8",
x"A5E17D91",
x"A4327C36",
x"A2927AED",
x"A12879C7",
x"A01B78DD",
x"9F8D783E",
x"9F9277FC",
x"A035781D",
x"A169789C",
x"A310796B",
x"A4FB7A74",
x"A6FA7B98",
x"A8D17CB7",
x"AA4D7DB0",
x"AB457E6A",
x"ABA17ED1",
x"AB5C7EDE",
x"AA847E95",
x"A9357E05",
x"A7997D41",
x"A5DE7C65",
x"A4327B8B",
x"A2BB7AC9",
x"A1977A33",
x"A0D779D4",
x"A08479B2",
x"A09A79CA",
x"A10B7A15",
x"A1C87A88",
x"A2B97B15",
x"A3C77BAD",
x"A4E07C41",
x"A5EB7CC6",
x"A6D97D30",
x"A79C7D7A",
x"A82E7D9F",
x"A8887DA0",
x"A8AF7D82",
x"A8A97D4E",
x"A8857D0F",
x"A8507CD0",
x"A81B7C9E",
x"A7F47C85",
x"A7EB7C8F",
x"A8077CC1",
x"A8497D1F",
x"A8AC7DA2",
x"A9297E46",
x"A9B27EFE",
x"AA397FBF",
x"AAAF807A",
x"AB0A8121",
x"AB4281A5",
x"AB568200",
x"AB498229",
x"AB218222",
x"AAE781ED",
x"AAA88195",
x"AA6B8126",
x"AA3B80B0",
x"AA188040",
x"AA057FE7",
x"A9FD7FAB",
x"A9F37F8F",
x"A9DA7F8E",
x"A9A57F9F",
x"A9437FAD",
x"A8AB7FAB",
x"A7D37F7F",
x"A6BA7F1F",
x"A5677E82",
x"A3E47DA5",
x"A2437C8F",
x"A0947B51",
x"9EE779FC",
x"9D4878A0",
x"9BB3774B",
x"9A247603",
x"988374C3",
x"96B3737C",
x"9495721D",
x"9205708D",
x"8EED6EB7",
x"8B3E6C8D",
x"86FC6A10",
x"82416748",
x"7D3A6455",
x"7824615C",
x"73475E8E",
x"6EE95C21",
x"6B525A3D",
x"68B5590C",
x"6733589E",
x"66D658F5",
x"67915A02",
x"69415BA4",
x"6BAE5DAB",
x"6E9B5FE7",
x"71C76224",
x"74F26435",
x"77E865F7",
x"7A806755",
x"7CA56848",
x"7E4B68D8",
x"7F756916",
x"8031691A",
x"80966901",
x"80BC68E5",
x"80BE68D9",
x"80B568EB",
x"80B76921",
x"80D56979",
x"811B69EC",
x"81916A6C",
x"82386AEF",
x"830B6B6B",
x"84036BD9",
x"85116C37",
x"86286C84",
x"87376CC5",
x"882F6D00",
x"89046D35",
x"89A96D66",
x"8A1A6D92",
x"8A536DB3",
x"8A586DC4",
x"8A2C6DBF",
x"89DC6DA1",
x"89706D6C",
x"88F66D26",
x"88776CD7",
x"87FE6C8C",
x"87966C54",
x"87426C3A",
x"87066C45",
x"86E56C76",
x"86D96CC7",
x"86E06D27",
x"86F36D86",
x"87076DCE",
x"87146DEF",
x"870E6DD8",
x"86ED6D86",
x"86A86CF9",
x"863B6C3D",
x"85A46B62",
x"84E76A80",
x"840B69AA",
x"831E68F6",
x"822B6873",
x"8146682B",
x"80816820",
x"7FEF684E",
x"7F9D68B0",
x"7F986938",
x"7FE769DE",
x"808A6A96",
x"817D6B59",
x"82B56C1E",
x"84216CE6",
x"85B16DAD",
x"874D6E72",
x"88E96F35",
x"8A6F6FF8",
x"8BD670B9",
x"8D187175",
x"8E327229",
x"8F2872D1",
x"8FFD7365",
x"90B673DF",
x"91597439",
x"91E47467",
x"92587461",
x"92AB7425",
x"92D673AC",
x"92CF72F9",
x"928D720F",
x"920A70F9",
x"91496FC8",
x"90506E8C",
x"8F2E6D5C",
x"8DF46C4F",
x"8CB96B78",
x"8B946AE5",
x"8A986A9E",
x"89D26AA8",
x"89466AFA",
x"88F36B83",
x"88CC6C31",
x"88C16CE9",
x"88B96D93",
x"88A56E17",
x"88726E65",
x"88146E6F",
x"87886E34",
x"86D36DB8",
x"86006D06",
x"85206C2E",
x"84426B48",
x"837C6A65",
x"82D9699A",
x"826868F7",
x"822A6886",
x"821D6849",
x"82396841",
x"82726862",
x"82B4689B",
x"82EA68DC",
x"8300690C",
x"82DC6914",
x"826A68E1",
x"819D6862",
x"8065678E",
x"7EC16666",
x"7CB564F3",
x"7A536348",
x"77B1617E",
x"74F25FB7",
x"723A5E12",
x"6FB25CB2",
x"6D835BB1",
x"6BCC5B1C",
x"6AAA5AFE",
x"6A2B5B50",
x"6A555C04",
x"6B215CFE",
x"6C7F5E27",
x"6E585F60",
x"70916093",
x"730D61AE",
x"75AE62AD",
x"785B6390",
x"7AFA6465",
x"7D76653A",
x"7FC16620",
x"81C86725",
x"83876852",
x"84F669A4",
x"86146B13",
x"86EA6C8A",
x"87806DF5",
x"87E76F38",
x"88347040",
x"887A70FC",
x"88CF7166",
x"89457185",
x"89E77162",
x"8ABF7113",
x"8BC570AE",
x"8CF3704E",
x"8E367003",
x"8F7C6FDB",
x"90AE6FD9",
x"91B86FFE",
x"928D703E",
x"93227090",
x"937A70E8",
x"939A713B",
x"93927186",
x"937671C8",
x"935A7209",
x"9356724D",
x"937A729D",
x"93D672FF",
x"94717376",
x"954C7400",
x"9660749A",
x"97A7753B",
x"991575DB",
x"9A9E7672",
x"9C3976FE",
x"9DDF777E",
x"9F8877F5",
x"A1327868",
x"A2D678DD",
x"A470795A",
x"A5F479DE",
x"A75A7A6A",
x"A8947AF5",
x"A9957B77",
x"AA547BEA",
x"AACF7C44",
x"AB077C86",
x"AB0A7CB3",
x"AAED7CD4",
x"AAD17CFA",
x"AAD77D36",
x"AB227D9F",
x"ABD27E4A",
x"AD027F43",
x"AEC2809B",
x"B118824F",
x"B3FE845D",
x"B76786B8",
x"BB39894F",
x"BF578C08",
x"C39F8ECE",
x"C7F09182",
x"CC23940A",
x"D0189651",
x"D3AA9841",
x"D6BD99CB",
x"D9349AE4",
x"DAF69B8A",
x"DBF69BBD",
x"DC299B86",
x"DB8B9AEE",
x"DA249A05",
x"D80898D8",
x"D54B9778",
x"D21395F3",
x"CE849456",
x"CACA92AE",
x"C713910A",
x"C38F8F77",
x"C0688E04",
x"BDC38CC2",
x"BBC08BC0",
x"BA6E8B10",
x"B9D68AB6",
x"B9EA8AB8",
x"BA958B0B",
x"BBAD8BA1",
x"BD028C59",
x"BE5B8D13",
x"BF7F8DA4",
x"C03D8DEC",
x"C06A8DC9",
x"BFF08D2F",
x"BECB8C1D",
x"BD0C8AA1",
x"BAD188D8",
x"B84586EA",
x"B5958500",
x"B2F0833F",
x"B07581C3",
x"AE388096",
x"AC357FB3",
x"AA517EFF",
x"A8677E57",
x"A6437D88",
x"A3AB7C67",
x"A0707AC9",
x"9C6C7896",
x"978E75C4",
x"91E07261",
x"8B896E88",
x"84BF6A6B",
x"7DD6663F",
x"77256245",
x"71075EB5",
x"6BCC5BC0",
x"67B5598B",
x"64E95828",
x"6376579B",
x"635157D7",
x"645458C3",
x"664C5A40",
x"68FF5C28",
x"6C2E5E55",
x"6FA760A7",
x"733B6300",
x"76D1654B",
x"7A556779",
x"7DC46982",
x"811E6B61",
x"84666D17",
x"879E6EA4",
x"8AC17009",
x"8DC5714A",
x"909E7264",
x"933C735B",
x"9590742F",
x"978B74E2",
x"99297578",
x"9A6B75F6",
x"9B5A7667",
x"9C0776D0",
x"9C82773C",
x"9CE677B0",
x"9D467836",
x"9DB878CD",
x"9E487975",
x"9EFB7A28",
x"9FD67AD7",
x"A0CA7B79",
x"A1CD7BFE",
x"A2C57C54",
x"A3987C71",
x"A42E7C4A",
x"A46C7BDE",
x"A43F7B33",
x"A39F7A54",
x"A2907953",
x"A11E7847",
x"9F69774A",
x"9D957675",
x"9BD275DA",
x"9A497586",
x"99247581",
x"987B75C1",
x"985A763A",
x"98BB76D4",
x"997E7774",
x"9A7D77FE",
x"9B877854",
x"9C647867",
x"9CE77826",
x"9CED7792",
x"9C6476B3",
x"9B4C759C",
x"99B97461",
x"97CD7321",
x"95B271F5",
x"939770F6",
x"91A77033",
x"90066FB7",
x"8ECB6F83",
x"8E006F92",
x"8DA76FD5",
x"8DB47043",
x"8E1770C8",
x"8EBF715A",
x"8F9871EE",
x"90977280",
x"91AF730F",
x"92DA739D",
x"94157431",
x"956274D2",
x"96BB758B",
x"9822765B",
x"9991774B",
x"9B037858",
x"9C6C797E",
x"9DC27AAF",
x"9EFA7BE0",
x"A0057CFC",
x"A0DF7DF1",
x"A17B7EAA",
x"A1D77F15",
x"A1F87F29",
x"A1E17EE3",
x"A19E7E43",
x"A13F7D5E",
x"A0DA7C4C",
x"A0817B2F",
x"A04C7A29",
x"A04C7960",
x"A08E78F1",
x"A11A78EE",
x"A1ED7960",
x"A2FE7A3A",
x"A43D7B6B",
x"A5927CD0",
x"A6E67E44",
x"A81E7F9F",
x"A92880C5",
x"A9F38199",
x"AA778214",
x"AAB38236",
x"AAB2820F",
x"AA8081B2",
x"AA298139",
x"A9C080BC",
x"A951804A",
x"A8E47FED",
x"A8777FA0",
x"A8007F59",
x"A76D7F02",
x"A6A47E85",
x"A5847DC6",
x"A3EE7CB3",
x"A1C67B3C",
x"9EF77960",
x"9B747723",
x"97487497",
x"928471D4",
x"8D536EF9",
x"87E96C28",
x"82846980",
x"7D6C671E",
x"78E0651B",
x"751E638A",
x"72536273",
x"709A61D8",
x"6FFC61B5",
x"706D6200",
x"71D162A8",
x"73FC639E",
x"76BA64CC",
x"79D56621",
x"7D1B678A",
x"805C68F9",
x"83776A61",
x"86526BBA",
x"88DF6D00",
x"8B1D6E33",
x"8D106F52",
x"8EC57062",
x"904B7166",
x"91AF725F",
x"92FE7351",
x"943F7437",
x"9570750D",
x"968E75D0",
x"978E7674",
x"986376F5",
x"98FE7750",
x"99597783",
x"99707793",
x"9948778C",
x"98F1777C",
x"98887772",
x"982B7781",
x"97FD77B3",
x"98187810",
x"98957898",
x"99797941",
x"9ABC79F9",
x"9C457AAC",
x"9DF37B43",
x"9F997BAD",
x"A1157BDE",
x"A2437BD9",
x"A3157BA6",
x"A38A7B60",
x"A3B57B20",
x"A3B87B0C",
x"A3BC7B3E",
x"A3EE7BD0",
x"A4747CC9",
x"A5667E28",
x"A6CD7FDD",
x"A89E81D1",
x"AAC283E4",
x"AD1285F3",
x"AF6487DF",
x"B192898E",
x"B37B8AF4",
x"B5078C06",
x"B6298CC5",
x"B6E38D34",
x"B73F8D5D",
x"B74C8D48",
x"B71F8D01",
x"B6D08C94",
x"B6758C10",
x"B6298B88",
x"B6028B14",
x"B6188ACC",
x"B67F8AC8",
x"B7468B1E",
x"B8748BDD",
x"BA028D06",
x"BBE18E8B",
x"BDF29052",
x"C00B9232",
x"C1FB93FA",
x"C391957A",
x"C4A09687",
x"C50E9706",
x"C4D196EB",
x"C3F5963F",
x"C29B9521",
x"C0EE93B7",
x"BF289231",
x"BD7790B7",
x"BC048F69",
x"BAE48E56",
x"BA188D7B",
x"B9898CC3",
x"B9168C0E",
x"B8958B3B",
x"B7DE8A29",
x"B6D788CC",
x"B5778721",
x"B3CD853F",
x"B1F8834A",
x"B02B8174",
x"AE987FF1",
x"AD747EF1",
x"ACE67E91",
x"ACFA7EDE",
x"ADA67FD0",
x"AECD8147",
x"B03A8314",
x"B1AD84FA",
x"B2E786BF",
x"B3AD882B",
x"B3DC8918",
x"B361896D",
x"B2468927",
x"B0A88853",
x"AEB3870E",
x"AC9E857E",
x"AA9283C6",
x"A8B3820B",
x"A7118061",
x"A59E7ED4",
x"A4387D5E",
x"A2A87BEB",
x"A0AB7A60",
x"9DFB7899",
x"9A607678",
x"95B573E4",
x"8FF370D2",
x"89356D47",
x"81BC695C",
x"79E3653B",
x"721D611A",
x"6AE15D3B",
x"64A359D9",
x"5FC5572F",
x"5C8A5566",
x"5B115491",
x"5B5154AD",
x"5D1E55A6",
x"602E574F",
x"64275971",
x"68A65BD5",
x"6D4E5E3D",
x"71D16081",
x"75F3627D",
x"79946421",
x"7CA4656D",
x"7F2A666F",
x"81356738",
x"82DE67E3",
x"843B6883",
x"855F6928",
x"865669DB",
x"87256A99",
x"87CC6B5E",
x"88496C1D",
x"889A6CCD",
x"88C16D62",
x"88C36DD5",
x"88AD6E24",
x"888D6E4F",
x"88736E5B",
x"88726E4B",
x"88916E29",
x"88D86DF8",
x"89436DBD",
x"89CC6D7F",
x"8A606D3F",
x"8AEF6D03",
x"8B656CCD",
x"8BAE6C9E",
x"8BC06C79",
x"8B976C5F",
x"8B356C51",
x"8AA56C4D",
x"89F96C51",
x"89426C5C",
x"88976C69",
x"88076C78",
x"879E6C84",
x"87606C8D",
x"87496C94",
x"874F6C94",
x"87606C90",
x"876D6C82",
x"87666C68",
x"873E6C3E",
x"86ED6C02",
x"86776BB2",
x"85E36B54",
x"853E6AE5",
x"84956A72",
x"83FA6A00",
x"8377699A",
x"83146947",
x"82CF690C",
x"82A368EC",
x"828068E2",
x"825968E8",
x"822068F5",
x"81C368FC",
x"813E68F6",
x"808E68DC",
x"7FBA68AB",
x"7ECE6863",
x"7DDF680D",
x"7D0167AE",
x"7C4C674F",
x"7BD366F9",
x"7BA166B1",
x"7BBC6679",
x"7C216650",
x"7CC46634",
x"7D8D6620",
x"7E676611",
x"7F376604",
x"7FE065F9",
x"804F65F0",
x"807465EC",
x"804965F2",
x"7FD265FF",
x"7F1D6614",
x"7E3C6630",
x"7D4C6649",
x"7C65665B",
x"7BA0665E",
x"7B13664B",
x"7ACE6621",
x"7AD365E6",
x"7B25659E",
x"7BBB6556",
x"7C87651E",
x"7D7C6503",
x"7E876511",
x"7F9A654F",
x"80A865BF",
x"81A8665B",
x"82916717",
x"836067E0",
x"841068A7",
x"84A06958",
x"850D69E2",
x"85596A3E",
x"85816A66",
x"858B6A5E",
x"85776A2B",
x"854869D9",
x"85016973",
x"84A768FF",
x"84346884",
x"83A56803",
x"82F06776",
x"820766D3",
x"80DB6613",
x"7F586527",
x"7D756407",
x"7B2A62AF",
x"787D6122",
x"757F5F6C",
x"724F5D9B",
x"6F175BC9",
x"6C075A12",
x"69545895",
x"672A576D",
x"65B056B0",
x"64FC5670",
x"651656B0",
x"65EE576E",
x"6769589B",
x"695F5A24",
x"6BA05BEA",
x"6DFD5DCF",
x"704A5FB3",
x"7266617D",
x"743E6313",
x"75C56468",
x"77036573",
x"78046635",
x"78DB66B8",
x"799D6706",
x"7A5D6731",
x"7B2B6749",
x"7C0E6762",
x"7D096786",
x"7E1467C2",
x"7F27681D",
x"8037689B",
x"8135693C",
x"821B69FC",
x"82E26AD5",
x"83896BBD",
x"84186CAD",
x"849A6D99",
x"851D6E76",
x"85AE6F3B",
x"865D6FDF",
x"87327058",
x"883270A0",
x"895970B4",
x"8A9E7093",
x"8BF4703E",
x"8D486FBE",
x"8E876F1D",
x"8FA26E69",
x"908E6DB3",
x"91436D0C",
x"91C26C84",
x"92116C2E",
x"92386C13",
x"92406C35",
x"92386C97",
x"92276D30",
x"92106DF3",
x"91FA6ED1",
x"91E26FB5",
x"91C97090",
x"91AC7152",
x"918A71F0",
x"91647265",
x"913B72B3",
x"910E72DC",
x"90E272EA",
x"90B572E1",
x"908A72CA",
x"905C72AB",
x"902B7285",
x"8FF37257",
x"8FB2721C",
x"8F6A71D1",
x"8F1E7174",
x"8ECF7103",
x"8E877082",
x"8E4D6FF8",
x"8E2B6F72",
x"8E276EFE",
x"8E456EA9",
x"8E8A6E80",
x"8EF36E8F",
x"8F7C6ED5",
x"901D6F52",
x"90CF6FF9",
x"918570BD",
x"92397186",
x"92E07243",
x"937372DE",
x"93EC7348",
x"94497379",
x"948B7374",
x"94B2733D",
x"94C272E6",
x"94BE7282",
x"94A77226",
x"948071E4",
x"944871CA",
x"93FB71DE",
x"9398721D",
x"931A727C",
x"927D72EA",
x"91C37352",
x"90F173A1",
x"900E73CA",
x"8F2773C4",
x"8E4C738D",
x"8D8E7333",
x"8CF972C3",
x"8C977251",
x"8C6971F4",
x"8C6C71BD",
x"8C8E71B9",
x"8CC171E8",
x"8CED7248",
x"8CFE72CB",
x"8CE7735E",
x"8C9E73EB",
x"8C25745F",
x"8B8474A9",
x"8ACB74BB",
x"8A097492",
x"894E742D",
x"889D7390",
x"87F272C3",
x"873E71C8",
x"866570A9",
x"85446F64",
x"83BB6DFC",
x"81AE6C6F",
x"7F0B6ABB",
x"7BD968E6",
x"782D66F7",
x"743764FC",
x"70326309",
x"6C6D6137",
x"69315FA5",
x"66C55E6D",
x"655C5DA7",
x"65165D63",
x"65F65DA8",
x"67E65E71",
x"6ABA5FAF",
x"6E306148",
x"7202631D",
x"75E9650A",
x"79A866F0",
x"7D0D68B1",
x"7FF96A38",
x"82606B79",
x"84496C72",
x"85C66D27",
x"86F36DA7",
x"87EC6E02",
x"88D06E47",
x"89B86E88",
x"8AB46ED2",
x"8BCE6F30",
x"8D066FA4",
x"8E59702B",
x"8FBF70C1",
x"9129715B",
x"928D71EB",
x"93D97266",
x"950372C3",
x"960172F8",
x"96CB7302",
x"975F72E2",
x"97BF72A1",
x"97F1724B",
x"980071EE",
x"97F7719C",
x"97E77164",
x"97DD7154",
x"97E67172",
x"980A71C3",
x"984C723E",
x"98AB72DC",
x"991F738B",
x"99A27437",
x"9A2674CE",
x"9A9F7541",
x"9B017582",
x"9B45758C",
x"9B647560",
x"9B607503",
x"9B3B7486",
x"9AF973F8",
x"9AA5736E",
x"9A4A72FF",
x"99F472BE",
x"99AE72BD",
x"99817306",
x"9976739D",
x"998E7480",
x"99CA75A2",
x"9A2676EE",
x"9A98784A",
x"9B117999",
x"9B817ABA",
x"9BD77B95",
x"9C077C12",
x"9C047C28",
x"9BCB7BD6",
x"9B5C7B29",
x"9AC07A3A",
x"9A0B7923",
x"994D7808",
x"989F7706",
x"98177639",
x"97C375B3",
x"97B17579",
x"97DF7589",
x"984575D4",
x"98D37646",
x"996F76C7",
x"99FA773E",
x"9A57779B",
x"9A6F77CD",
x"9A2B77CE",
x"9985779F",
x"98837744",
x"973276CB",
x"95AE763E",
x"941A75AC",
x"9297751F",
x"914B74A1",
x"904F743A",
x"8FB873EE",
x"8F8A73BD",
x"8FC373A9",
x"905573B1",
x"912873D4",
x"92297412",
x"93407468",
x"946074D7",
x"957D755B",
x"969475EF",
x"97A97690",
x"98BE7733",
x"99D677CD",
x"9AED7851",
x"9BF878AF",
x"9CE978DB",
x"9DA578CA",
x"9E177875",
x"9E2577DB",
x"9DC37703",
x"9CEC75FB",
x"9BA974D5",
x"9A1073AA",
x"983B728D",
x"96497195",
x"945770CA",
x"92797033",
x"90B16FC4",
x"8EF76F6C",
x"8D346F12",
x"8B466E94",
x"890D6DD8",
x"866A6CC5",
x"83506B4F",
x"7FC46977",
x"7BDB674E",
x"77C664F0",
x"73C16286",
x"7010603C",
x"6CF65E41",
x"6AAA5CB9",
x"69525BBF",
x"68FD5B61",
x"69A35B9E",
x"6B275C64",
x"6D5E5D9C",
x"70145F27",
x"731760E2",
x"763E62B1",
x"7968647D",
x"7C866638",
x"7F9467DB",
x"82976968",
x"859A6AE3",
x"88A76C57",
x"8BC26DC7",
x"8EEA6F3A",
x"921570B0",
x"95317226",
x"98297396",
x"9AE774F6",
x"9D577640",
x"9F71776C",
x"A12E7874",
x"A2927958",
x"A3AB7A18",
x"A48B7ABA",
x"A5487B43",
x"A5F87BBA",
x"A6B07C29",
x"A77F7C96",
x"A8737D09",
x"A98B7D85",
x"AAC77E0F",
x"AC1F7EAA",
x"AD847F56",
x"AEEA8012",
x"B03F80D9",
x"B17081A8",
x"B2728276",
x"B33D833B",
x"B3D283EE",
x"B432848A",
x"B46D8505",
x"B495855C",
x"B4C0858D",
x"B5048598",
x"B5738585",
x"B618855C",
x"B6F58527",
x"B80784F1",
x"B93A84C7",
x"BA7884B3",
x"BBA584BD",
x"BCA284E6",
x"BD57852B",
x"BDAC8582",
x"BD9485E2",
x"BD098635",
x"BC13866E",
x"BABC867A",
x"B918864C",
x"B74085E2",
x"B554853B",
x"B3748463",
x"B1C28370",
x"B0608278",
x"AF6D8198",
x"AEFF80EB",
x"AF288085",
x"AFEB8075",
x"B13F80BF",
x"B30B8159",
x"B5298230",
x"B768832D",
x"B9928432",
x"BB6E851E",
x"BCC985D6",
x"BD7E8646",
x"BD77865E",
x"BCB4861B",
x"BB468581",
x"B94F849B",
x"B6FA8378",
x"B47A8230",
x"B1FC80D3",
x"AFA67F77",
x"AD917E2A",
x"ABC67CFA",
x"AA407BED",
x"A8F47B08",
x"A7CC7A4D",
x"A6B579B6",
x"A59E793E",
x"A47E78E1",
x"A3537896",
x"A2247857",
x"A0F9781F",
x"9FDF77EA",
x"9EE077B3",
x"9E03777C",
x"9D437744",
x"9C9A7708",
x"9BFA76C7",
x"9B507682",
x"9A917634",
x"99AE75E0",
x"989F7581",
x"976C7519",
x"961A74AC",
x"94BC743D",
x"936673D1",
x"922C736F",
x"911E731A",
x"904572D5",
x"8FA2729C",
x"8F2C726A",
x"8ECD7230",
x"8E6971E2",
x"8DDB716B",
x"8CFE70BB",
x"8BB16FC3",
x"89D66E78",
x"875F6CD8",
x"84496AEC",
x"80A468C2",
x"7C916673",
x"783F6418",
x"73E661D5",
x"6FCA5FC6",
x"6C265E08",
x"69345CB2",
x"67235BD2",
x"660D5B6D",
x"65F95B81",
x"66D95C06",
x"68905CE9",
x"6AEF5E17",
x"6DBD5F77",
x"70C160F6",
x"73C46279",
x"769763ED",
x"791D6546",
x"7B416677",
x"7D03677C",
x"7E6D6854",
x"7F906904",
x"80866997",
x"81656A16",
x"82416A8A",
x"83286AFD",
x"84216B76",
x"852A6BF6",
x"863C6C7C",
x"874B6D00",
x"884C6D7A",
x"89356DE3",
x"89FD6E30",
x"8AA26E5E",
x"8B256E6C",
x"8B896E61",
x"8BD56E44",
x"8C0D6E26",
x"8C386E13",
x"8C586E17",
x"8C6F6E3A",
x"8C7D6E7D",
x"8C816EDB",
x"8C7B6F4A",
x"8C6D6FB7",
x"8C5A7013",
x"8C48704B",
x"8C3E7055",
x"8C45702B",
x"8C636FD2",
x"8C9E6F57",
x"8CF66EC7",
x"8D676E3B",
x"8DE96DC8",
x"8E6F6D7F",
x"8EEA6D69",
x"8F4F6D8C",
x"8F8E6DDF",
x"8FA26E54",
x"8F846ED5",
x"8F396F4D",
x"8EC66FA4",
x"8E386FC7",
x"8D9A6FAB",
x"8CFB6F4E",
x"8C6D6EB3",
x"8BF76DE6",
x"8BA56CFF",
x"8B7D6C12",
x"8B7D6B37",
x"8BA56A87",
x"8BEF6A13",
x"8C4F69E5",
x"8CBB6A00",
x"8D256A63",
x"8D806B00",
x"8DBE6BC7",
x"8DD66CA1",
x"8DC26D7C",
x"8D7E6E43",
x"8D106EE2",
x"8C7D6F54",
x"8BD26F90",
x"8B1B6F9A",
x"8A6A6F7A",
x"89C96F3B",
x"89426EEC",
x"88DA6E9A",
x"88906E4E",
x"885C6E12",
x"88326DE6",
x"88066DCD",
x"87C66DC1",
x"87696DBA",
x"86E66DB3",
x"86396DA1",
x"85656D82",
x"84736D4E",
x"836D6D04",
x"82656CA7",
x"81656C34",
x"80796BB0",
x"7FAA6B1D",
x"7EF96A7F",
x"7E6269D9",
x"7DDF6931",
x"7D686889",
x"7CED67E5",
x"7C6A674B",
x"7BD866BF",
x"7B326646",
x"7A7E65E3",
x"79C46598",
x"79096566",
x"785C6548",
x"77C6653C",
x"774E653B",
x"76F7653E",
x"76BE653E",
x"769A652F",
x"767F650E",
x"765864CF",
x"7613646D",
x"759963E2",
x"74D86327",
x"73BD6237",
x"723D610E",
x"704F5FAE",
x"6DF65E1A",
x"6B3B5C57",
x"68315A76",
x"64F35888",
x"61A356A4",
x"5E6C54E7",
x"5B7D536B",
x"5903524D",
x"572A51A0",
x"56125174",
x"55D151C9",
x"566B5295",
x"57D553C4",
x"59EE5538",
x"5C8956C7",
x"5F6F584D",
x"626259A2",
x"65285AA9",
x"67905B52",
x"69795B95",
x"6ACE5B80",
x"6B935B25",
x"6BD75AA4",
x"6BBA5A1E",
x"6B6159B5",
x"6AF25984",
x"6A8F5998",
x"6A5259F6",
x"6A4C5A95",
x"6A7D5B64",
x"6AE35C48",
x"6B705D27",
x"6C145DE6",
x"6CBE5E73",
x"6D635EC5",
x"6DFA5ED7",
x"6E805EAF",
x"6EF35E5A",
x"6F585DE4",
x"6FB45D5F",
x"70095CD5",
x"705B5C50",
x"70AB5BDA",
x"70F65B77",
x"713B5B29",
x"71775AF6",
x"71A85AE0",
x"71CC5AEB",
x"71E65B1E",
x"71F65B78",
x"72005BFD",
x"72065CA7",
x"720C5D71",
x"72145E4F",
x"72205F35",
x"72306011",
x"724560D9",
x"72616181",
x"72826206",
x"72AA6266",
x"72DB62A7",
x"731762D2",
x"735F62F0",
x"73B26309",
x"74116321",
x"74796338",
x"74E26349",
x"7548634E",
x"75A3633B",
x"75E9630B",
x"761662B8",
x"76256245",
x"761461B7",
x"75E6611B",
x"759E6084",
x"75486006",
x"74EA5FB1",
x"74945F95",
x"744E5FBB",
x"74216022",
x"741760C5",
x"74316198",
x"74726289",
x"74D56384",
x"75546474",
x"75E8654B",
x"768765F9",
x"772B6676",
x"77C966BE",
x"786066D5",
x"78E966BE",
x"79636683",
x"79D1662E",
x"7A3165C8",
x"7A8A655E",
x"7ADC64F7",
x"7B2A64A0",
x"7B74645A",
x"7BBC642F",
x"7C04641E",
x"7C496427",
x"7C8E6449",
x"7CD26480",
x"7D1A64C5",
x"7D686514",
x"7DC16568",
x"7E2B65BA",
x"7EAB6609",
x"7F446652",
x"7FF66696",
x"80BE66D3",
x"8197670E",
x"82736746",
x"8346677A",
x"840167AA",
x"849467D1",
x"84F467ED",
x"851867FA",
x"850067F5",
x"84B167DE",
x"843867B4",
x"83A2677C",
x"83016738",
x"826566F0",
x"81D566A5",
x"8152665B",
x"80D3660B",
x"804465B5",
x"7F8A654E",
x"7E8764C8",
x"7D1E641B",
x"7B39633B",
x"78D16224",
x"75E860D6",
x"72975F5C",
x"6F045DC1",
x"6B635C1B",
x"67EF5A85",
x"64E1591A",
x"626B57EE",
x"60B15718",
x"5FCA56A1",
x"5FB1568B",
x"605656D3",
x"61935767",
x"633B5838",
x"651E592C",
x"670D5A2E",
x"68E15B2B",
x"6A825C14",
x"6BE15CE0",
x"6CFD5D8B",
x"6DE55E1A",
x"6EA85E8E",
x"6F585EF1",
x"70065F49",
x"70BE5F9D",
x"71845FED",
x"7255603C",
x"73276088",
x"73ED60D0",
x"749B6113",
x"7524614F",
x"75806183",
x"75AE61B4",
x"75B261E3",
x"759A6217",
x"756F624F",
x"75446291",
x"752762DA",
x"7521632D",
x"753C6383",
x"757A63D8",
x"75D66428",
x"764C646C",
x"76D264A0",
x"775F64BF",
x"77ED64CB",
x"787964C1",
x"790164A5",
x"79896480",
x"7A106455",
x"7A9D642F",
x"7B32641A",
x"7BCF641E",
x"7C706444",
x"7D106491",
x"7DA7650A",
x"7E2E65AB",
x"7EA16670",
x"7EFF674E",
x"7F486835",
x"7F846917",
x"7FC169E5",
x"80096A90",
x"80696B10",
x"80E96B61",
x"818D6B84",
x"82536B83",
x"83326B66",
x"841B6B3B",
x"84FA6B0D",
x"85BC6AE8",
x"86506ACF",
x"86AC6AC8",
x"86C96AD2",
x"86AC6AE8",
x"86656B07",
x"86036B2A",
x"85A06B4F",
x"85526B75",
x"85326B9C",
x"854F6BC7",
x"85B56BF6",
x"86656C2D",
x"87586C68",
x"887E6CA6",
x"89C66CE1",
x"8B186D16",
x"8C5F6D3F",
x"8D846D5E",
x"8E776D6C",
x"8F2C6D6F",
x"8F9E6D68",
x"8FCB6D5B",
x"8FB86D4B",
x"8F6A6D38",
x"8EEF6D20",
x"8E4F6D00",
x"8D976CD1",
x"8CD36C8F",
x"8C0D6C35",
x"8B4E6BC7",
x"8A9D6B47",
x"8A016AC2",
x"89846A47",
x"892569E3",
x"88EC69A7",
x"88D969A0",
x"88EA69D1",
x"891F6A37",
x"896F6AC7",
x"89D26B70",
x"8A396C1C",
x"8A9A6CB1",
x"8AE36D19",
x"8B066D41",
x"8AF76D21",
x"8AAF6CB8",
x"8A2F6C0F",
x"897C6B32",
x"889E6A38",
x"87A76935",
x"86A5683F",
x"85AA6763",
x"84BB66A8",
x"83DC6610",
x"83016590",
x"821A651A",
x"81076495",
x"7FAA63F0",
x"7DDF6313",
x"7B8D61EF",
x"78A6607A",
x"752A5EB8",
x"71305CB5",
x"6CDE5A87",
x"686B584D",
x"6419562C",
x"602B5447",
x"5CE152C2",
x"5A6C51B7",
x"58E95139",
x"5864514A",
x"58CA51E1",
x"59F952EB",
x"5BC15447",
x"5DE655D3",
x"602B5767",
x"625C58E1",
x"644D5A28",
x"65DF5B26",
x"67075BD5",
x"67C55C35",
x"68275C53",
x"68405C3D",
x"682A5C0A",
x"67FD5BCC",
x"67D25B91",
x"67BB5B67",
x"67C55B56",
x"67F55B5D",
x"684E5B7B",
x"68CC5BA9",
x"69695BE3",
x"6A1C5C1F",
x"6AD85C57",
x"6B935C87",
x"6C425CA9",
x"6CDE5CC2",
x"6D625CCD",
x"6DCF5CD2",
x"6E275CD3",
x"6E735CD9",
x"6EBE5CEC",
x"6F165D12",
x"6F855D56",
x"70165DBD",
x"70CC5E4D",
x"71AA5F04",
x"72A85FDF",
x"73BA60D5",
x"74CF61D8",
x"75D662D8",
x"76BE63C5",
x"7776648B",
x"77F3651E",
x"78346573",
x"783A6587",
x"7810655C",
x"77C464FD",
x"77686477",
x"770D63DF",
x"76C86346",
x"76A462C4",
x"76AD6266",
x"76E3623C",
x"7749624C",
x"77D36294",
x"787A630D",
x"792D63AB",
x"79DD645C",
x"7A80650D",
x"7B0765A7",
x"7B6C661A",
x"7BAE6658",
x"7BCE6659",
x"7BD26620",
x"7BC565B4",
x"7BAF6525",
x"7B9B6489",
x"7B9063F9",
x"7B8C6389",
x"7B90634F",
x"7B936356",
x"7B8E63A3",
x"7B76642D",
x"7B4564E3",
x"7AF465B1",
x"7A8A667D",
x"7A0C672D",
x"798A67AB",
x"791767E9",
x"78C567E5",
x"78A867A0",
x"78CB672B",
x"79316697",
x"79D865FD",
x"7AB16570",
x"7BA56503",
x"7C9E64BE",
x"7D7D64A4",
x"7E2864AF",
x"7E8E64D5",
x"7EA0650A",
x"7E5F653C",
x"7DD06562",
x"7D096573",
x"7C1A656C",
x"7B21654F",
x"7A346523",
x"796964ED",
x"78CF64BB",
x"786D6490",
x"78416473",
x"78426465",
x"78656463",
x"7898646A",
x"78CC6474",
x"78F3647D",
x"7901647F",
x"78F06476",
x"78BC6465",
x"78696446",
x"77F96420",
x"776D63ED",
x"76C863AD",
x"760A635A",
x"753162F4",
x"743D6273",
x"732B61D3",
x"72026115",
x"70C8603E",
x"6F8C5F58",
x"6E625E71",
x"6D655D9F",
x"6CAD5CF7",
x"6C535C8D",
x"6C6C5C74",
x"6CFF5CB6",
x"6E0D5D57",
x"6F8C5E50",
x"71655F91",
x"737F6106",
x"75BB6293",
x"77FF6423",
x"7A3765A1",
x"7C566703",
x"7E5F6842",
x"805F6968",
x"826A6A7D",
x"849A6B96",
x"87086CC5",
x"89C96E1A",
x"8CE76FA1",
x"9062715B",
x"94267344",
x"981A754B",
x"9C157760",
x"9FED7965",
x"A3747B47",
x"A6837CED",
x"A8FD7E47",
x"AAD67F4D",
x"AC127FFE",
x"ACC78064",
x"AD18808C",
x"AD35808E",
x"AD568082",
x"ADAC8081",
x"AE6780A5",
x"AFA980FE",
x"B180819B",
x"B3E7827D",
x"B6C7839F",
x"B9FB84F4",
x"BD4E8666",
x"C08787DD",
x"C3728942",
x"C5E58A7B",
x"C7C48B7D",
x"C9088C3E",
x"C9B98CC1",
x"C9F78D0D",
x"C9EA8D36",
x"C9C48D52",
x"C9B68D73",
x"C9EA8DAC",
x"CA798E07",
x"CB728E8A",
x"CCCD8F2E",
x"CE748FE9",
x"D04090AA",
x"D2099162",
x"D3A39200",
x"D4E49279",
x"D5AA92C7",
x"D5E892E8",
x"D59692E0",
x"D4BE92B9",
x"D376927C",
x"D1DE922F",
x"D01891DD",
x"CE4A918E",
x"CC9A9144",
x"CB299101",
x"CA0E90CB",
x"C95890A0",
x"C9129084",
x"C9369077",
x"C9B9907A",
x"CA86908A",
x"CB7F90A5",
x"CC8490C7",
x"CD7190E2",
x"CE2390ED",
x"CE7F90E0",
x"CE6C90AE",
x"CDDD904E",
x"CCD08FBB",
x"CB4A8EF4",
x"C95A8DFE",
x"C7158CDD",
x"C4918B9B",
x"C1E78A42",
x"BF2988DF",
x"BC678778",
x"B9A98618",
x"B6F384C5",
x"B4438380",
x"B199824A",
x"AEF58123",
x"AC5A8008",
x"A9C97EF5",
x"A7527DE4",
x"A5017CD6",
x"A2E77BC7",
x"A1147ABA",
x"9F9479B7",
x"9E7078C3",
x"9DA977E8",
x"9D397731",
x"9D1476A9",
x"9D257652",
x"9D577633",
x"9D917646",
x"9DB9767F",
x"9DBD76D2",
x"9D90772A",
x"9D287777",
x"9C8A77A5",
x"9BBB77A9",
x"9ACC7781",
x"99CF772F",
x"98D676BD",
x"97ED7639",
x"971D75B1",
x"965D752F",
x"959F74B4",
x"94C3743D",
x"93A573B9",
x"9215730C",
x"8FED721F",
x"8D0A70D2",
x"89586F16",
x"84DC6CE1",
x"7FAF6A3A",
x"7A036737",
x"742163FF",
x"6E5C60C2",
x"69105DB6",
x"64935B0D",
x"613058F1",
x"5F175781",
x"5E6356C7",
x"5F0F56C0",
x"60F6575A",
x"63E55875",
x"679059EB",
x"6BA85B95",
x"6FE05D53",
x"73EF5F07",
x"779D609D",
x"7AC2620D",
x"7D486352",
x"7F2A6470",
x"8073656C",
x"8138664B",
x"81966710",
x"81A867BC",
x"81916851",
x"816868C8",
x"81436921",
x"8134695B",
x"813F6973",
x"81686972",
x"81A7695B",
x"81F46938",
x"82456914",
x"828B68F9",
x"82BE68EC",
x"82D568F3",
x"82D06911",
x"82B46942",
x"82876980",
x"825569C2",
x"822D69FF",
x"82156A2D",
x"821A6A44",
x"82396A3F",
x"82706A20",
x"82B869E8",
x"8303699D",
x"8345694B",
x"837668FC",
x"839168BE",
x"839A689B",
x"839B68A1",
x"83A268D2",
x"83C56931",
x"841569BC",
x"84A26A6C",
x"85766B37",
x"868D6C0D",
x"87DF6CE5",
x"89596DB1",
x"8AE36E66",
x"8C5D6F00",
x"8DAE6F7C",
x"8EBC6FDB",
x"8F767024",
x"8FD0705F",
x"8FCB7093",
x"8F6C70C7",
x"8EC570FF",
x"8DE6713A",
x"8CE97176",
x"8BE571AF",
x"8AF171DA",
x"8A2471EF",
x"898E71E9",
x"893C71C3",
x"89397179",
x"89837112",
x"8A147090",
x"8AE06FFC",
x"8BD66F5F",
x"8CDF6EC4",
x"8DE26E31",
x"8EC66DAE",
x"8F796D41",
x"8FEC6CEE",
x"90186CB7",
x"90046C9D",
x"8FBB6CA1",
x"8F536CC4",
x"8EE46D04",
x"8E876D5E",
x"8E526DCD",
x"8E536E47",
x"8E916EC5",
x"8F066F40",
x"8FA46FA9",
x"90596FFC",
x"910B7034",
x"91A77054",
x"921B705F",
x"92627061",
x"927A7064",
x"926F7073",
x"9252709C",
x"923670E1",
x"92327143",
x"924F71B9",
x"92937234",
x"92F672A0",
x"936972E6",
x"93D372F2",
x"941A72B1",
x"9420721C",
x"93D07133",
x"93217002",
x"92106E9C",
x"90A86D1D",
x"8EFD6BA4",
x"8D256A4E",
x"8B3E6932",
x"8959685F",
x"878767D6",
x"85CC6791",
x"8424677A",
x"82846779",
x"80DF6770",
x"7F2A6744",
x"7D5E66DE",
x"7B7C6635",
x"79936549",
x"77BA642B",
x"760B62EF",
x"74A761B4",
x"73A8609D",
x"73275FC8",
x"73305F4D",
x"73C15F3E",
x"74D25F9B",
x"76526060",
x"782A617E",
x"7A3F62DF",
x"7C80646C",
x"7EDC6610",
x"814C67B7",
x"83CF6955",
x"866C6AE8",
x"89296C6B",
x"8C106DE5",
x"8F246F5C",
x"926470D5",
x"95C97254",
x"994673DA",
x"9CC57565",
x"A02E76EF",
x"A3697871",
x"A66079E3",
x"A9057B3D",
x"AB4F7C7C",
x"AD3D7D9E",
x"AEDE7EA2",
x"B0407F8B",
x"B17B8061",
x"B2A88129",
x"B3DA81E8",
x"B52282A5",
x"B68A835C",
x"B80E840E",
x"B9A284B3",
x"BB338546",
x"BCA385BD",
x"BDD7860F",
x"BEB58635",
x"BF23862C",
x"BF1985F3",
x"BE988592",
x"BDA98515",
x"BC65848D",
x"BAF08408",
x"B970839E",
x"B80B835D",
x"B6E88353",
x"B6288384",
x"B5DD83F1",
x"B6148494",
x"B6C9855A",
x"B7F28636",
x"B9788711",
x"BB4287D6",
x"BD298877",
x"BF1188E4",
x"C0D38917",
x"C254890E",
x"C37B88CC",
x"C4338859",
x"C47787C0",
x"C444870F",
x"C3A68657",
x"C2AF85A5",
x"C17B850D",
x"C02C849E",
x"BEE78467",
x"BDD18476",
x"BD0884D0",
x"BCA3857B",
x"BCB28673",
x"BD3087AC",
x"BE118914",
x"BF3A8A93",
x"C08B8C0D",
x"C1DD8D66",
x"C3088E83",
x"C3EF8F4C",
x"C47C8FB7",
x"C4A28FB9",
x"C4638F5B",
x"C3CC8EA5",
x"C2EF8DAC",
x"C1E88C84",
x"C0CE8B46",
x"BFB68A07",
x"BEAF88D8",
x"BDBC87C6",
x"BCDE86D9",
x"BC0C8614",
x"BB3A8576",
x"BA5E84FA",
x"B96E849C",
x"B867845A",
x"B74F842F",
x"B62F8417",
x"B5198411",
x"B425841C",
x"B3678439",
x"B2F28463",
x"B2D4849B",
x"B31184DD",
x"B3A38523",
x"B47B8568",
x"B57F85A2",
x"B68B85C9",
x"B77A85D4",
x"B82385BC",
x"B8688578",
x"B82F850A",
x"B768846E",
x"B61683AB",
x"B44782C5",
x"B21281C5",
x"AF9580B3",
x"ACEE7F95",
x"AA327E6D",
x"A76E7D35",
x"A4A17BE5",
x"A1B67A72",
x"9E9278CD",
x"9B0E76E7",
x"970774B4",
x"92637230",
x"8D1D6F61",
x"87416C54",
x"80FA6923",
x"7A8765EF",
x"743B62E0",
x"6E6A601F",
x"696D5DCF",
x"65895C0E",
x"62EC5AF1",
x"61A65A7B",
x"61AA5AA6",
x"62CC5B5D",
x"64CE5C82",
x"67645DF1",
x"6A3B5F84",
x"6D116118",
x"6FAD628E",
x"71E863D2",
x"73AF64D5",
x"75066598",
x"75F96620",
x"769E6675",
x"771466A8",
x"777066C8",
x"77C966E2",
x"782E66FF",
x"78A86724",
x"793B6756",
x"79E66791",
x"7AA767D5",
x"7B79681B",
x"7C566860",
x"7D3868A0",
x"7E1768D6",
x"7EEB6900",
x"7FA86919",
x"8046691E",
x"80BC690C",
x"810468E2",
x"811D68A0",
x"81076848",
x"80D167E0",
x"80866775",
x"803B6711",
x"800466C5",
x"7FF766A0",
x"802166AD",
x"808966F2",
x"812F676D",
x"820A6817",
x"830768DF",
x"840E69B1",
x"85066A76",
x"85D26B19",
x"86636B8A",
x"86AC6BC2",
x"86AF6BC4",
x"86776B97",
x"86186B51",
x"85AE6B04",
x"85536ACB",
x"85226AB7",
x"852E6AD2",
x"857A6B20",
x"86046B9C",
x"86BB6C34",
x"87876CD8",
x"884C6D70",
x"88EF6DE9",
x"895A6E34",
x"89836E47",
x"896A6E21",
x"891A6DCB",
x"88AB6D54",
x"88356CCB",
x"87D86C45",
x"87AA6BD7",
x"87BF6B8F",
x"88206B79",
x"88C66BA0",
x"89AD6C04",
x"8ABC6CA6",
x"8BE36D7D",
x"8D086E83",
x"8E1C6FA9",
x"8F0D70E1",
x"8FD27219",
x"90667341",
x"90C97446",
x"90FA7516",
x"90FB75A2",
x"90CE75DE",
x"907075C6",
x"8FE37554",
x"8F277490",
x"8E3B7385",
x"8D24723E",
x"8BE670D2",
x"8A8B6F54",
x"89226DD8",
x"87B76C6D",
x"86586B27",
x"85186A10",
x"8403692E",
x"83276887",
x"828D6820",
x"823867F6",
x"822D680C",
x"8262685C",
x"82D368E6",
x"837069A4",
x"842A6A8C",
x"84E96B90",
x"859D6CA1",
x"86316DAD",
x"86966E9E",
x"86C26F62",
x"86B46FE6",
x"86697020",
x"85EC7009",
x"85426FA1",
x"84766EEF",
x"838B6DFC",
x"82816CD4",
x"814F6B82",
x"7FE66A0D",
x"7E35687A",
x"7C2566C6",
x"79AA64F2",
x"76BA62F7",
x"735B60D9",
x"6FA55E9B",
x"6BBD5C4F",
x"67D55A07",
x"642857E6",
x"60F65609",
x"5E795496",
x"5CDF53A9",
x"5C475354",
x"5CBA53A2",
x"5E2E5487",
x"608555ED",
x"638F57B6",
x"671459B9",
x"6AD75BCD",
x"6E9D5DCF",
x"72375FA5",
x"757D6141",
x"785962A1",
x"7AC463CE",
x"7CBF64D6",
x"7E5C65D0",
x"7FAE66C9",
x"80CE67CE",
x"81D268DC",
x"82CB69EF",
x"83C56AF7",
x"84C56BDF",
x"85C86C92",
x"86C66D00",
x"87B26D1E",
x"887D6CEC",
x"891B6C72",
x"89806BBF",
x"89A56AEC",
x"898B6A11",
x"89376945",
x"88AF689B",
x"88066826",
x"874867E9",
x"868367E6",
x"85C46819",
x"85136877",
x"847468F9",
x"83E56991",
x"83626A35",
x"82E36ADC",
x"82606B7D",
x"81D26C10",
x"81356C90",
x"80896CF5",
x"7FCF6D38",
x"7F136D59",
x"7E5B6D54",
x"7DB46D27",
x"7D2A6CD7",
x"7CC66C68",
x"7C906BE3",
x"7C8A6B52",
x"7CB16ABF",
x"7CFD6A35",
x"7D6569BA",
x"7DD86952",
x"7E466901",
x"7E9E68C2",
x"7ED36894",
x"7EDB686F",
x"7EB0684E",
x"7E566827",
x"7DD667F9",
x"7D3E67BE",
x"7C9D6775",
x"7C00671A",
x"7B7766AD",
x"7B06662E",
x"7AAE659E",
x"7A6564FD",
x"7A236452",
x"79D963A1",
x"798062F3",
x"79136259",
x"789D61E0",
x"7830619B",
x"77EB619E",
x"77EF61F4",
x"786562AB",
x"796A63C1",
x"7B166531",
x"7D6A66EB",
x"805C68D8",
x"83C96ADB",
x"87876CD7",
x"8B5C6EAE",
x"8F127051",
x"927971B0",
x"956D72CB",
x"97DA73AC",
x"99BF7461",
x"9B257501",
x"9C24759D",
x"9CD67647",
x"9D557705",
x"9DB177D5",
x"9DF478A9",
x"9E1B796D",
x"9E1E7A06",
x"9DEC7A5E",
x"9D767A5E",
x"9CB379FB",
x"9BA17936",
x"9A467819",
x"98B476BC",
x"9701753D",
x"954C73BE",
x"93B27261",
x"92507141",
x"91397075",
x"907C7005",
x"901B6FF0",
x"90117031",
x"904F70B5",
x"90BC7166",
x"913F722B",
x"91B272EB",
x"91EF738B",
x"91D073F2",
x"9132740C",
x"8FF473C7",
x"8E007313",
x"8B4C71EB",
x"87DD704E",
x"83CB6E47",
x"7F3E6BE9",
x"7A6F6952",
x"759D66A5",
x"7113640B",
x"6D1361AF",
x"69D65FB8",
x"67895E3F",
x"663F5D59",
x"65F65D07",
x"66975D41",
x"67F85DEC",
x"69E35EE9",
x"6C236017",
x"6E7D614E",
x"70C76272",
x"72DF636A",
x"74B5642F",
x"764864BC",
x"77A0651B",
x"78CF6559",
x"79EA6584",
x"7B0465AF",
x"7C2B65E9",
x"7D686638",
x"7EBA66A4",
x"801E672D",
x"818B67D1",
x"82F46889",
x"844F694E",
x"858E6A17",
x"86AC6ADC",
x"87A46B94",
x"886F6C33",
x"890E6CB1",
x"89816D06",
x"89C96D2A",
x"89E66D1A",
x"89D96CD8",
x"89A56C63",
x"894E6BC8",
x"88D56B13",
x"88426A54",
x"879D699C",
x"86EF68FD",
x"86426886",
x"85A06844",
x"8514683B",
x"84A8686C",
x"846268D1",
x"8446695F",
x"84556A0C",
x"848E6AC5",
x"84EA6B82",
x"85636C33",
x"85F16CD2",
x"868E6D5F",
x"87356DD8",
x"87E66E41",
x"88A16EA4",
x"896C6F06",
x"8A4F6F6E",
x"8B4E6FDE",
x"8C6D7057",
x"8DAA70D5",
x"8EFC7152",
x"905871C7",
x"91A8722A",
x"92D97274",
x"93D7729F",
x"949072AB",
x"94FA729C",
x"9517727B",
x"94F07250",
x"94977227",
x"9425720C",
x"93B57205",
x"935D7216",
x"932F723E",
x"93347278",
x"936672BA",
x"93B872FB",
x"94177330",
x"946A7352",
x"9497735E",
x"948A7354",
x"94387339",
x"939A7312",
x"92B972E8",
x"91A172BE",
x"90647299",
x"8F187274",
x"8DD27248",
x"8CA1720F",
x"8B9371BE",
x"8AAE714F",
x"89F670BE",
x"89687012",
x"89016F52",
x"88BC6E93",
x"88916DE6",
x"887C6D61",
x"88746D14",
x"88736D09",
x"88726D3F",
x"88696DAD",
x"88526E3E",
x"88256ED4",
x"87DF6F52",
x"877D6F9A",
x"87016F96",
x"86716F34",
x"85D36E78",
x"852F6D6B",
x"84936C26",
x"84046AC8",
x"838B6976",
x"832A6854",
x"82E0677C",
x"82A86701",
x"827966E8",
x"82456724",
x"81FD67A0",
x"81906838",
x"80EC68C5",
x"7FFF691D",
x"7EBB6919",
x"7D19689E",
x"7B13679E",
x"78AD661B",
x"75F36424",
x"72FC61D8",
x"6FE25F60",
x"6CCB5CED",
x"69DF5AAF",
x"674558D2",
x"65275774",
x"63A056AC",
x"62C85681",
x"62A856E7",
x"633E57CC",
x"6478590E",
x"663D5A8B",
x"686C5C21",
x"6AE15DAF",
x"6D755F1A",
x"700A6055",
x"72866158",
x"74DB6225",
x"76FD62CB",
x"78F26356",
x"7ABD63D8",
x"7C696465",
x"7E016507",
x"7F9065CC",
x"811866B8",
x"829D67C9",
x"841868F9",
x"85836A3D",
x"86D16B87",
x"87FA6CCA",
x"88F46DF6",
x"89BF6F00",
x"8A596FDE",
x"8AC9708A",
x"8B1E7105",
x"8B657151",
x"8BAE7175",
x"8C097179",
x"8C7E7166",
x"8D127145",
x"8DC1711F",
x"8E7D70F8",
x"8F3870D4",
x"8FDC70B4",
x"90537097",
x"908B707F",
x"90797065",
x"9018704B",
x"8F6E702D",
x"8E88700D",
x"8D7D6FE9",
x"8C656FC3",
x"8B5A6F94",
x"8A776F61",
x"89CC6F24",
x"89646EDE",
x"89426E8A",
x"895F6E2D",
x"89AD6DC5",
x"8A186D58",
x"8A8E6CEE",
x"8AFB6C8C",
x"8B4E6C3B",
x"8B7A6C04",
x"8B776BE9",
x"8B466BEF",
x"8AE76C10",
x"8A646C47",
x"89C86C89",
x"891E6CCA",
x"88746CFC",
x"87D96D14",
x"875B6D09",
x"87066CD8",
x"86E56C80",
x"86FE6C09",
x"87596B7D",
x"87F26AE9",
x"88C36A5E",
x"89C269E9",
x"8ADD6994",
x"8BFE696B",
x"8D0D696C",
x"8DF46996",
x"8EA169E2",
x"8F066A47",
x"8F1D6ABA",
x"8EED6B2E",
x"8E866B9E",
x"8DFA6C03",
x"8D666C5F",
x"8CE56CB5",
x"8C8D6D0C",
x"8C6D6D69",
x"8C8D6DD5",
x"8CE36E52",
x"8D606EDE",
x"8DEA6F76",
x"8E63700D",
x"8EAB7097",
x"8EAF7106",
x"8E62714D",
x"8DC57164",
x"8CEA7145",
x"8BED70F6",
x"8AF67080",
x"8A286FEE",
x"89A86F51",
x"898D6EBA",
x"89E36E35",
x"8A9F6DCD",
x"8BAC6D86",
x"8CE76D61",
x"8E246D59",
x"8F3C6D6B",
x"900B6D8F",
x"90806DBF",
x"90936DFA",
x"904D6E3E",
x"8FC36E89",
x"8F106ED7",
x"8E4B6F23",
x"8D816F66",
x"8CB96F92",
x"8BE56F96",
x"8AEA6F5E",
x"89A26ED8",
x"87E96DF3",
x"859B6CA8",
x"82A56AF3",
x"7F0368DF",
x"7AC9667C",
x"762163E6",
x"7145613E",
x"6C795EA7",
x"68055C46",
x"64275A38",
x"61145897",
x"5EEE5771",
x"5DC056CC",
x"5D8656A6",
x"5E2956F1",
x"5F87579E",
x"617C5891",
x"63DF59B6",
x"66875AF1",
x"69565C2C",
x"6C2E5D55",
x"6EF75E5C",
x"719E5F3C",
x"74135FF2",
x"764A6084",
x"783C60FE",
x"79E66170",
x"7B4C61E9",
x"7C77627D",
x"7D7A633E",
x"7E6C6432",
x"7F626563",
x"807966CC",
x"81C16863",
x"83486A17",
x"850B6BD1",
x"87016D76",
x"89116EF0",
x"8B1A7029",
x"8CF9710F",
x"8E87719A",
x"8FA771CD",
x"904371AD",
x"9058714B",
x"8FE970BA",
x"8F0E7010",
x"8DE56F5F",
x"8C906EB8",
x"8B326E29",
x"89EC6DB1",
x"88D56D54",
x"87F76D0A",
x"87586CCD",
x"86F06C93",
x"86B46C57",
x"86916C12",
x"867D6BC2",
x"866A6B6B",
x"86536B0F",
x"86356AB5",
x"86136A62",
x"85F06A1C",
x"85D669E5",
x"85C869C1",
x"85C869B0",
x"85D569B0",
x"85ED69C1",
x"860B69DF",
x"862C6A0A",
x"864B6A3F",
x"86656A7D",
x"867C6AC1",
x"86946B09",
x"86B76B51",
x"86E96B99",
x"87346BDE",
x"879E6C21",
x"882B6C62",
x"88DF6CA4",
x"89B76CEB",
x"8AAF6D3B",
x"8BC46D9C",
x"8CEF6E12",
x"8E2A6EA0",
x"8F6D6F4A",
x"90B4700D",
x"91F670E8",
x"932C71D2",
x"945272C5",
x"955D73B7",
x"9646749A",
x"97067565",
x"9792760D",
x"97E67688",
x"97FE76CE",
x"97DA76DD",
x"977B76B3",
x"96E97652",
x"962C75C7",
x"9550751A",
x"9465745E",
x"937373A3",
x"928A72FB",
x"91B27275",
x"90F3721C",
x"905071F5",
x"8FCC71FF",
x"8F647231",
x"8F1A727B",
x"8EE972CB",
x"8ECF730D",
x"8EC97331",
x"8ED57329",
x"8EEC72EC",
x"8F0A727C",
x"8F2771E1",
x"8F387126",
x"8F34705C",
x"8F0E6F96",
x"8EBE6EE5",
x"8E3B6E57",
x"8D836DEF",
x"8C976DB0",
x"8B7A6D92",
x"8A356D8A",
x"88CE6D85",
x"874B6D70",
x"85AC6D37",
x"83F26CC8",
x"82116C16",
x"80006B17",
x"7DB469C9",
x"7B236832",
x"7846665F",
x"7528645D",
x"71D56245",
x"6E68602B",
x"6B045E28",
x"67D45C4D",
x"64FD5AAE",
x"62A65950",
x"60E85839",
x"5FD45769",
x"5F6856D6",
x"5F975678",
x"604A5646",
x"61595632",
x"62A75635",
x"640F564C",
x"65735673",
x"66BF56AF",
x"67EC5704",
x"68F75777",
x"69E6580B",
x"6AC858C3",
x"6BA6599E",
x"6C8C5A97",
x"6D835BA4",
x"6E895CB8",
x"6F9B5DC9",
x"70B05EC8",
x"71B55FA9",
x"72A06064",
x"736060F6",
x"73ED615A",
x"74426195",
x"746261AE",
x"745261A8",
x"7425618E",
x"73EA6168",
x"73B8613B",
x"73A0610B",
x"73B160DC",
x"73F360B1",
x"74686088",
x"750A6064",
x"75CB6045",
x"7699602B",
x"775E6018",
x"7804600E",
x"787C6010",
x"78B8601E",
x"78B5603C",
x"78796069",
x"780D60A4",
x"778460E9",
x"76F66139",
x"76756191",
x"761361EC",
x"75DF624B",
x"75DF62AB",
x"7610630E",
x"76696374",
x"76DC63DF",
x"7752644C",
x"77BA64B8",
x"77FF651E",
x"78146576",
x"77F065B8",
x"779665DC",
x"770965DB",
x"765865AE",
x"75946556",
x"74D464D9",
x"7427643E",
x"73A06394",
x"734562EA",
x"731D6250",
x"732461D5",
x"734E6183",
x"738E6160",
x"73D66170",
x"741961AE",
x"74496213",
x"74656293",
x"746A6323",
x"746063B7",
x"744F6444",
x"744264C2",
x"74446527",
x"745B656F",
x"74876595",
x"74C46594",
x"7509656D",
x"7547651E",
x"757064A8",
x"75756410",
x"754C635F",
x"74F3629B",
x"746961D2",
x"73B8610E",
x"72EF605A",
x"721E5FBE",
x"71595F3E",
x"70B05EDA",
x"702B5E92",
x"6FD55E5D",
x"6FAB5E35",
x"6FA75E10",
x"6FBE5DE7",
x"6FDF5DB6",
x"6FFC5D7A",
x"70035D31",
x"6FE55CDD",
x"6F995C82",
x"6F195C22",
x"6E655BBF",
x"6D845B5A",
x"6C825AF4",
x"6B6B5A8E",
x"6A545A29",
x"694C59C6",
x"68635969",
x"67A75915",
x"671A58CD",
x"66BD5894",
x"66845867",
x"66615843",
x"663B581F",
x"65FA57F0",
x"658457A8",
x"64C4573A",
x"63A8569C",
x"622B55CA",
x"605554C4",
x"5E345396",
x"5BE95250",
x"5997510B",
x"57694FE2",
x"558C4EF4",
x"54264E57",
x"53584E1F",
x"53374E56",
x"53CA4EFC",
x"5509500B",
x"56E2516D",
x"5935530C",
x"5BDC54CE",
x"5EAE5699",
x"61835852",
x"643759E6",
x"66AA5B45",
x"68CB5C67",
x"6A8F5D49",
x"6BF25DEE",
x"6CF95E5D",
x"6DAF5E9D",
x"6E235EB8",
x"6E605EB7",
x"6E7A5EA1",
x"6E7C5E80",
x"6E755E5A",
x"6E725E33",
x"6E7A5E0E",
x"6E9A5DED",
x"6ED45DD0",
x"6F2D5DB8",
x"6FA45DA4",
x"70375D94",
x"70DB5D87",
x"71895D7D",
x"72345D7A",
x"72CF5D80",
x"73525D92",
x"73B55DB6",
x"73F35DF0",
x"740E5E41",
x"74075EAB",
x"73E55F2B",
x"73AB5FBC",
x"735F6056",
x"730460EC",
x"729D6174",
x"722661E0",
x"719E6228",
x"710A6245",
x"70696237",
x"6FC46200",
x"6F2561AE",
x"6E9E614E",
x"6E3D60F2",
x"6E1160A8",
x"6E2A6083",
x"6E8A608B",
x"6F3460C3",
x"70196129",
x"712861B1",
x"72496248",
x"736062D9",
x"744F634F",
x"75026397",
x"7563639E",
x"75706360",
x"752D62DD",
x"74A4621E",
x"73ED6137",
x"7327603C",
x"726C5F4C",
x"71DB5E7E",
x"718A5DEA",
x"71895DA1",
x"71DD5DA9",
x"72865E04",
x"73725EA4",
x"748D5F78",
x"75BC606C",
x"76E36163",
x"77E86248",
x"78B06306",
x"79286390",
x"794B63DF",
x"791463F6",
x"788A63DA",
x"77BC639B",
x"76BE6345",
x"75A362E4",
x"74826286",
x"736F622F",
x"727D61E6",
x"71B761A5",
x"7123616A",
x"70C4612E",
x"709660EE",
x"709160A7",
x"70AE6058",
x"70E26007",
x"71215FB9",
x"71655F7C",
x"71A75F56",
x"71E35F55",
x"721A5F7C",
x"724C5FCF",
x"7280604F",
x"72B760F6",
x"72F761B9",
x"73426290",
x"739A6369",
x"73FD643B",
x"746964F6",
x"74DB6590",
x"754B6601",
x"75B56645",
x"76116655",
x"765B6632",
x"768765DF",
x"7690655E",
x"766964B4",
x"760963E8",
x"75636300",
x"74736201",
x"733260F6",
x"71A15FE2",
x"6FCB5ECF",
x"6DC15DC2",
x"6B9E5CC5",
x"69835BDF",
x"67975B18",
x"65FC5A7A",
x"64D25A0B",
x"643159D5",
x"642159D7",
x"64A05A17",
x"659D5A92",
x"66FF5B46",
x"68A75C2B",
x"6A775D36",
x"6C555E62",
x"6E305F9F",
x"700060E9",
x"71C96238",
x"739A6389",
x"758364D9",
x"7798662E",
x"79EC6789",
x"7C8968ED",
x"7F706A61",
x"829E6BE2",
x"86046D6F",
x"89906F02",
x"8D277092",
x"90B27213",
x"9418737E",
x"974374C3",
x"9A1E75DE",
x"9C9A76C7",
x"9EAE7782",
x"A052780F",
x"A188787B",
x"A25678CE",
x"A2C97919",
x"A2F37964",
x"A2E979BC",
x"A2C67A26",
x"A2A47AA3",
x"A2977B30",
x"A2B17BC4",
x"A2FB7C56",
x"A3787CD7",
x"A4217D40",
x"A4EA7D85",
x"A5C37DA6",
x"A6987DA2",
x"A7597D7F",
x"A7F87D49",
x"A86E7D08",
x"A8B87CC9",
x"A8D77C95",
x"A8D07C6F",
x"A8AE7C5E",
x"A8757C5B",
x"A8327C64",
x"A7E97C74",
x"A79F7C84",
x"A7597C92",
x"A7147C9C",
x"A6CF7CA0",
x"A6877CA2",
x"A6327C9C",
x"A5C87C8F",
x"A53B7C77",
x"A4827C4D",
x"A3947C09",
x"A26B7BA3",
x"A1077B16",
x"9F717A63",
x"9DB5798B",
x"9BE97896",
x"9A247793",
x"98807692",
x"971175A2",
x"95E774D0",
x"95067425",
x"946A73A3",
x"94077348",
x"93C97310",
x"939E72F1",
x"937072DF",
x"933672D8",
x"92EC72D7",
x"929472DF",
x"923F72F6",
x"91FB7321",
x"91E07366",
x"91F773C8",
x"924C7444",
x"92D974D0",
x"9394755C",
x"946775DB",
x"95367639",
x"95E77664",
x"96627654",
x"96947606",
x"96787581",
x"961474D0",
x"9577740C",
x"94B67348",
x"93F072A0",
x"933F7224",
x"92BB71E4",
x"927771E2",
x"927B721A",
x"92C67280",
x"934F7300",
x"94017385",
x"94C673F2",
x"95867436",
x"9622743E",
x"96887402",
x"96A5737E",
x"966E72B9",
x"95E271C1",
x"950470A9",
x"93E16F86",
x"928A6E6F",
x"91106D79",
x"8F836CB1",
x"8DED6C1E",
x"8C566BBE",
x"8AB66B83",
x"89016B59",
x"87206B21",
x"84F96ABB",
x"826F6A03",
x"7F6A68DC",
x"7BDF6735",
x"77C86504",
x"73386255",
x"6E4F5F41",
x"693E5BEE",
x"64425895",
x"5F9F5570",
x"5B9652B6",
x"5861509D",
x"562E4F4D",
x"55154ED7",
x"55194F3D",
x"5626506D",
x"58165242",
x"5AB6548C",
x"5DC55718",
x"610C59AF",
x"644F5C24",
x"67645E52",
x"6A2A6021",
x"6C936187",
x"6E9B6289",
x"704E632F",
x"71B8638D",
x"72F063B7",
x"740663C1",
x"750763BE",
x"75FC63BB",
x"76E663C4",
x"77C263DD",
x"7887640D",
x"79306453",
x"79B264AF",
x"7A10651E",
x"7A47659D",
x"7A5B6625",
x"7A5566B2",
x"7A42673F",
x"7A2B67C8",
x"7A1B6845",
x"7A1B68B2",
x"7A31690D",
x"7A5C6954",
x"7A9B6984",
x"7AEC699E",
x"7B4769A1",
x"7BA7698E",
x"7C066966",
x"7C606927",
x"7CB268D5",
x"7CFF6873",
x"7D466804",
x"7D8E6790",
x"7DDD671E",
x"7E3766BA",
x"7E9E666C",
x"7F16663F",
x"7F9B6638",
x"8028665E",
x"80B866AD",
x"813F6723",
x"81B567B8",
x"820E685F",
x"8248690D",
x"825969B5",
x"82466A49",
x"82146AC2",
x"81C66B1C",
x"816C6B57",
x"810E6B75",
x"80B96B7F",
x"80766B7C",
x"804C6B72",
x"80446B69",
x"805B6B62",
x"80936B5F",
x"80E96B5B",
x"815B6B4F",
x"81E36B37",
x"827D6B0D",
x"83236ACC",
x"83CC6A76",
x"84716A0F",
x"8509699C",
x"85866927",
x"85DC68BB",
x"86036862",
x"85ED6820",
x"859567FA",
x"84FA67EF",
x"841E67F9",
x"830B680D",
x"81CF6823",
x"807C682D",
x"7F276820",
x"7DE867F6",
x"7CD067A8",
x"7BF3673B",
x"7B5866B0",
x"7B036611",
x"7AEF6569",
x"7B1464C5",
x"7B60642F",
x"7BC263B2",
x"7C276356",
x"7C7C631D",
x"7CB46303",
x"7CC26306",
x"7CA36318",
x"7C566331",
x"7BDE6344",
x"7B3F6345",
x"7A80632A",
x"79A462EA",
x"78B16287",
x"77A86200",
x"768B615A",
x"755E609D",
x"74215FD0",
x"72DB5F00",
x"71935E36",
x"70555D78",
x"6F2A5CCD",
x"6E1E5C38",
x"6D385BB9",
x"6C795B4D",
x"6BD95AF1",
x"6B4E5AA1",
x"6AC25A55",
x"6A1D5A05",
x"694259AC",
x"681E593F",
x"66A058B9",
x"64C25815",
x"628C5751",
x"6011566D",
x"5D75556E",
x"5ADC5460",
x"58765351",
x"566E5257",
x"54E55187",
x"53F950F4",
x"53B650B6",
x"541C50DA",
x"551D5166",
x"56A35254",
x"5889539B",
x"5AAE5522",
x"5CEC56CA",
x"5F215875",
x"61335A04",
x"630D5B5A",
x"64A35C66",
x"65F35D1F",
x"67035D8B",
x"67DC5DB8",
x"688C5DBD",
x"69245DB8",
x"69B45DC1",
x"6A4A5DED",
x"6AF05E4C",
x"6BAB5EE0",
x"6C7F5FA1",
x"6D62607E",
x"6E4E615F",
x"6F356229",
x"700D62C5",
x"70C46321",
x"71536331",
x"71B162F9",
x"71DC6283",
x"71D661E3",
x"71A76131",
x"715C6084",
x"71015FF7",
x"70A85F97",
x"70605F70",
x"70385F7E",
x"703B5FBC",
x"706D601D",
x"70D2608D",
x"716560FD",
x"721E615F",
x"72F361AD",
x"73D661E2",
x"74BA6203",
x"7593621B",
x"76586238",
x"77076262",
x"779E62A7",
x"7820630B",
x"78936390",
x"78FF642E",
x"796964DC",
x"79D8658B",
x"7A4B662A",
x"7AC566AA",
x"7B4166FF",
x"7BBC6723",
x"7C2F6713",
x"7C9966D5",
x"7CF46670",
x"7D4265F3",
x"7D83656D",
x"7DBE64ED",
x"7DF36481",
x"7E2B6437",
x"7E696413",
x"7EAE641D",
x"7EFA6456",
x"7F4F64BE",
x"7FA76550",
x"80006606",
x"805566D3",
x"80A267B0",
x"80E6688A",
x"81186954",
x"813869FD",
x"81416A7A",
x"812F6ABD",
x"81036AC2",
x"80B96A89",
x"80536A1A",
x"7FD66980",
x"7F4568D1",
x"7EAA681D",
x"7E0A677A",
x"7D7066F9",
x"7CE666A1",
x"7C706677",
x"7C146675",
x"7BD26690",
x"7BA866B5",
x"7B9466D8",
x"7B9166E8",
x"7B9866DB",
x"7BA566B0",
x"7BB1666C",
x"7BB86618",
x"7BB765C8",
x"7BA76589",
x"7B876566",
x"7B51656A",
x"7B026594",
x"7A9665DB",
x"7A0C6630",
x"79656680",
x"78A666BA",
x"77D666C8",
x"76FF669E",
x"762E6637",
x"756C6593",
x"74C464BB",
x"743863BE",
x"73C862AB",
x"736C6193",
x"73176083",
x"72B85F81",
x"723A5E94",
x"718D5DB9",
x"70A75CF0",
x"6F855C2F",
x"6E2A5B77",
x"6CA85AC5",
x"6B1A5A1C",
x"699C5982",
x"684E5901",
x"675158A1",
x"66BD586B",
x"66A05867",
x"66FD5897",
x"67D158F8",
x"69055985",
x"6A825A35",
x"6C2B5AFA",
x"6DE25BC9",
x"6F8F5C98",
x"71195D5C",
x"72755E0E",
x"739A5EAE",
x"74875F3C",
x"75425FBB",
x"75D26031",
x"763F60A7",
x"76966122",
x"76DF61AB",
x"77256246",
x"777262F7",
x"77CC63BE",
x"783B6495",
x"78BF6579",
x"795D665B",
x"7A11672E",
x"7AD567E6",
x"7BA16870",
x"7C6A68C2",
x"7D2768D2",
x"7DCE689E",
x"7E5C682B",
x"7ECF6784",
x"7F3266BF",
x"7F8E65F3",
x"7FF4653E",
x"807664BA",
x"8122647F",
x"820364A0",
x"831B6523",
x"84626604",
x"85C9673B",
x"873868AB",
x"88976A3B",
x"89CB6BC8",
x"8ABC6D31",
x"8B606E5C",
x"8BB16F35",
x"8BB86FB4",
x"8B876FD9",
x"8B356FB1",
x"8AE26F54",
x"8AA76EDB",
x"8A9A6E61",
x"8AC96E00",
x"8B386DCD",
x"8BDD6DCE",
x"8CAA6E09",
x"8D866E73",
x"8E566EFE",
x"8F046F92",
x"8F7C701A",
x"8FAF7085",
x"8FA170C0",
x"8F5870C1",
x"8EE3708A",
x"8E59701F",
x"8DD36F89",
x"8D696ED8",
x"8D286E1A",
x"8D1D6D62",
x"8D496CBE",
x"8DA46C3A",
x"8E226BE1",
x"8EAF6BB7",
x"8F3B6BC2",
x"8FB26C06",
x"900B6C7D",
x"903F6D24",
x"904F6DF2",
x"90456EDB",
x"902C6FCF",
x"901370C3",
x"900471A0",
x"900A725B",
x"902972E8",
x"905D7340",
x"909F7361",
x"90E37351",
x"91177316",
x"912F72BB",
x"911D724A",
x"90D671CB",
x"90597144",
x"8FA770B7",
x"8EC97020",
x"8DCC6F80",
x"8CC26ED2",
x"8BBE6E1A",
x"8AD36D5B",
x"8A176CA1",
x"89976BFD",
x"895D6B80",
x"89726B3E",
x"89CE6B45",
x"8A6A6B9E",
x"8B346C47",
x"8C136D34",
x"8CEF6E4D",
x"8DAC6F73",
x"8E317085",
x"8E67715E",
x"8E4571E5",
x"8DC17202",
x"8CE071AF",
x"8BAC70EC",
x"8A326FCA",
x"887E6E5B",
x"869E6CB5",
x"84946AEF",
x"825C6919",
x"7FEA673B",
x"7D2D6558",
x"7A11636A",
x"76846169",
x"72805F4D",
x"6E095D11",
x"69355AB9",
x"642A5852",
x"5F1D55EE",
x"5A5053A9",
x"560351A3",
x"52784FFB",
x"4FDF4ECA",
x"4E574E22",
x"4DE94E09",
x"4E864E7C",
x"50084F6A",
x"523750BD",
x"54D75254",
x"57A65412",
x"5A6B55D7",
x"5CFB5787",
x"5F38590A",
x"611D5A55",
x"62AE5B5C",
x"63FD5C1F",
x"65265CA4",
x"663F5CF3",
x"67655D1B",
x"68A15D28",
x"69FC5D2E",
x"6B705D39",
x"6CF25D57",
x"6E6F5D94",
x"6FD55DF4",
x"71135E78",
x"72185F1B",
x"72DE5FD5",
x"73626094",
x"73A7614E",
x"73B561EF",
x"7397626A",
x"735962B5",
x"730962C9",
x"72B162A8",
x"725F6256",
x"721861DD",
x"71E96150",
x"71D260C1",
x"71D96042",
x"72025FE9",
x"72495FC2",
x"72B25FD8",
x"733B602F",
x"73DE60C6",
x"749A6191",
x"7568627E",
x"7645637D",
x"772B6473",
x"7814654C",
x"78FC65F7",
x"79DD6669",
x"7AB4669A",
x"7B796690",
x"7C2B6658",
x"7CC66600",
x"7D48659D",
x"7DAF6542",
x"7DFA6501",
x"7E2864E2",
x"7E3A64E8",
x"7E2E650E",
x"7E036549",
x"7DB86589",
x"7D4B65BC",
x"7CB865D5",
x"7BFC65C5",
x"7B16658B",
x"7A076527",
x"78D5649E",
x"778663FF",
x"76276355",
x"74C562AD",
x"73736211",
x"72416188",
x"713B6115",
x"706C60B5",
x"6FD86063",
x"6F7D601B",
x"6F545FD8",
x"6F4B5F97",
x"6F555F59",
x"6F5F5F1F",
x"6F5C5EF0",
x"6F425ED0",
x"6F0F5EC2",
x"6EC25EC9",
x"6E685EE0",
x"6E0A5F04",
x"6DBB5F2C",
x"6D845F4F",
x"6D705F64",
x"6D825F64",
x"6DB55F4F",
x"6E035F22",
x"6E5B5EE4",
x"6EB15EA1",
x"6EF55E60",
x"6F1D5E31",
x"6F245E1A",
x"6F0F5E25",
x"6EE35E52",
x"6EB15EA1",
x"6E8A5F0B",
x"6E7F5F86",
x"6E9D6007",
x"6EEC6083",
x"6F6D60EE",
x"701A6142",
x"70E36176",
x"71B7618A",
x"727F617D",
x"73256153",
x"739A6111",
x"73D260BF",
x"73CB6062",
x"73846000",
x"730A5F9E",
x"72685F42",
x"71AA5EEA",
x"70DB5E92",
x"6FFD5E35",
x"6F105DC8",
x"6E0A5D3D",
x"6CDE5C8B",
x"6B795BA8",
x"69CC5A8B",
x"67CF5936",
x"658057B2",
x"62EC560E",
x"602E5464",
x"5D6C52D3",
x"5ADA517C",
x"58AB5081",
x"57164FFB",
x"56444FFF",
x"56585093",
x"575B51AF",
x"59455340",
x"5BF85525",
x"5F425739",
x"62E95952",
x"66AB5B4C",
x"6A475D06",
x"6D835E6C",
x"70385F74",
x"72516025",
x"73C8608A",
x"74AD60B8",
x"751B60C3",
x"753860C1",
x"752760BF",
x"750D60C5",
x"750260D2",
x"751160DD",
x"753E60DC",
x"757A60C3",
x"75B7608A",
x"75DE602D",
x"75D95FB2",
x"759E5F24",
x"75275E95",
x"747C5E1E",
x"73AE5DD2",
x"72D65DC6",
x"72165E06",
x"718A5E94",
x"714E5F6D",
x"71756083",
x"720661C2",
x"72FC6311",
x"74496459",
x"75D56581",
x"777F667A",
x"792A6737",
x"7AB567B2",
x"7C0D67F0",
x"7D2567FA",
x"7DFD67DC",
x"7EA067A8",
x"7F1E6770",
x"7F966746",
x"801E6738",
x"80D26753",
x"81BF679D",
x"82ED6817",
x"845368BC",
x"85E26982",
x"877C6A5C",
x"89016B3A",
x"8A526C0A",
x"8B556CBF",
x"8BF96D4D",
x"8C396DAE",
x"8C226DE3",
x"8BC86DF3",
x"8B4B6DE9",
x"8ACB6DD1",
x"8A696DBA",
x"8A396DB1",
x"8A466DBE",
x"8A8B6DE5",
x"8AF76E21",
x"8B6C6E6C",
x"8BC86EBA",
x"8BEC6EF8",
x"8BBB6F1A",
x"8B286F13",
x"8A346EDB",
x"88EA6E6F",
x"87676DD1",
x"85CC6D0A",
x"843F6C28",
x"82E06B3A",
x"81CB6A51",
x"810A697A",
x"80A468C4",
x"808A6837",
x"80AB67D3",
x"80EF679D",
x"81386789",
x"81706793",
x"818367AE",
x"816667D1",
x"811667F3",
x"8091680D",
x"7FE5681A",
x"7F186814",
x"7E3B67FD",
x"7D5867D5",
x"7C79679B",
x"7BA86753",
x"7AE866FA",
x"7A386694",
x"79986620",
x"790365A0",
x"78726514",
x"77DC6481",
x"773A63EF",
x"7689635F",
x"75C462DA",
x"74EA6268",
x"7402620A",
x"730E61C2",
x"7217618E",
x"71236168",
x"703A6145",
x"6F5C611B",
x"6E8A60DF",
x"6DC16081",
x"6CF65FFE",
x"6C205F4F",
x"6B375E74",
x"6A315D74",
x"690C5C59",
x"67C85B32",
x"66705A0E",
x"651058FE",
x"63BB5812",
x"62835757",
x"617C56D4",
x"60B75691",
x"6040568C",
x"601D56C3",
x"6051572C",
x"60D657C0",
x"61A65874",
x"62B6593D",
x"63FC5A11",
x"656E5AE9",
x"67035BBF",
x"68B55C94",
x"6A825D69",
x"6C635E41",
x"6E595F21",
x"705F6010",
x"72726110",
x"748C6222",
x"76A46348",
x"78B76477",
x"7AB965A8",
x"7CA866CF",
x"7E7F67DE",
x"803C68CB",
x"81E3698D",
x"83776A20",
x"85036A84",
x"868E6AC1",
x"88216AE1",
x"89C56AF3",
x"8B7F6B09",
x"8D4F6B34",
x"8F376B80",
x"91326BFA",
x"933C6CA8",
x"954D6D8D",
x"975F6EA4",
x"99696FE8",
x"9B66714F",
x"9D5272D1",
x"9F28745F",
x"A0E675EF",
x"A2857775",
x"A40778E7",
x"A5677A3A",
x"A6A87B68",
x"A7CC7C6B",
x"A8D77D40",
x"A9D37DE7",
x"AACA7E63",
x"ABC97EB9",
x"ACD97EF0",
x"AE017F0F",
x"AF467F1F",
x"B09F7F25",
x"B2027F25",
x"B35E7F1F",
x"B49C7F15",
x"B5AB7F07",
x"B6777EF8",
x"B6FB7EE7",
x"B7397EDD",
x"B73F7EE1",
x"B7237EFE",
x"B7077F3F",
x"B70B7FB0",
x"B74F8059",
x"B7EB8139",
x"B8EE824F",
x"BA57838E",
x"BC1C84EA",
x"BE23864F",
x"C05187AC",
x"C28288F3",
x"C4988A12",
x"C6778B08",
x"C80C8BD0",
x"C9508C6F",
x"CA408CE7",
x"CAE18D43",
x"CB3C8D87",
x"CB5B8DB5",
x"CB498DCB",
x"CB0C8DC6",
x"CAAC8DA1",
x"CA298D55",
x"C9858CDF",
x"C8C08C40",
x"C7DA8B7E",
x"C6D38A9F",
x"C5A989B2",
x"C46088C0",
x"C2F787DA",
x"C16E8707",
x"BFC9864D",
x"BE0E85AE",
x"BC428527",
x"BA6E84B1",
x"B8A38446",
x"B6F183E0",
x"B56D837E",
x"B42B831E",
x"B33D82C7",
x"B2B3827E",
x"B291824A",
x"B2D38233",
x"B36B823B",
x"B440825C",
x"B5328291",
x"B61882CD",
x"B6CC82FE",
x"B7298314",
x"B71182FE",
x"B67382B1",
x"B5448225",
x"B38B815A",
x"B1518057",
x"AEAB7F22",
x"ABAD7DC9",
x"A8697C51",
x"A4ED7AC4",
x"A1437922",
x"9D70776A",
x"99707597",
x"954573A6",
x"90F07195",
x"8C7A6F64",
x"87F76D21",
x"83836ADE",
x"7F4468B2",
x"7B6866BF",
x"78186523",
x"758363F6",
x"73C4634E",
x"72EF632F",
x"73076398",
x"74026476",
x"75C565B1",
x"7832672A",
x"7B2568C4",
x"7E776A63",
x"820B6BF6",
x"85C66D76",
x"89986EE4",
x"8D79704B",
x"916271BB",
x"9556734A",
x"99597506",
x"9D6E76FF",
x"A19B793A",
x"A5E37BB3",
x"AA477E63",
x"AECA8135",
x"B36A8419",
x"B82086F7",
x"BCE489B5",
x"C1A38C3E",
x"C6468E80",
x"CAB2906D",
x"CECB91FF",
x"D2759332",
x"D59B9411",
x"D83094A7",
x"DA349507",
x"DBB39549",
x"DCC39584",
x"DD7E95D1",
x"DE039641",
x"DE6F96DF",
x"DED097AD",
x"DF2E98A1",
x"DF8599AB",
x"DFC79AB1",
x"DFE49B9A",
x"DFCA9C4B",
x"DF6C9CB1",
x"DECD9CC1",
x"DDF59C7B",
x"DCFC9BEB",
x"DC009B26",
x"DB239A45",
x"DA859966",
x"DA3E98A3",
x"DA5B9810",
x"DADB97B5",
x"DBAC9793",
x"DCB197A0",
x"DDC797CB",
x"DEBE97FC",
x"DF729820",
x"DFBD9823",
x"DF8597F9",
x"DEBD97A0",
x"DD6A971D",
x"DB9C967C",
x"D96F95D2",
x"D7109534",
x"D4AF94B7",
x"D27B946A",
x"D0A5945C",
x"CF54948D",
x"CEA394FA",
x"CE999599",
x"CF2F9656",
x"D048971D",
x"D1BC97D6",
x"D351986E",
x"D4D398CB",
x"D60698E5",
x"D6C398B0",
x"D6E5982B",
x"D667975E",
x"D54D9652",
x"D3B49520",
x"D1C693D9",
x"CFB3929D",
x"CDB09182",
x"CBED909E",
x"CA8C9003",
x"C9A98FBB",
x"C9478FC2",
x"C95E9010",
x"C9D79090",
x"CA909127",
x"CB6891B9",
x"CC39922B",
x"CCE89266",
x"CD65925F",
x"CDAC9213",
x"CDC6918E",
x"CDC390E7",
x"CDC1903E",
x"CDDA8FB2",
x"CE238F63",
x"CEAC8F67",
x"CF748FC9",
x"D06E9087",
x"D17F918D",
x"D28992BF",
x"D36593F8",
x"D3F59510",
x"D42295E3",
x"D3E59659",
x"D3469666",
x"D2559607",
x"D132954C",
x"CFF49447",
x"CEB0930D",
x"CD6A91B5",
x"CC109048",
x"CA7E8EC6",
x"C87A8D22",
x"C5C48B46",
x"C21D8917",
x"BD51867A",
x"B749835E",
x"B00A7FC2",
x"A7C67BB3",
x"9ECA7754",
x"958B72D8",
x"8C876E7F",
x"84416A8A",
x"7D2E6738",
x"77AB64B7",
x"73EA6323",
x"71FC6280",
x"71BF62BC",
x"72FA63B2",
x"7554652D",
x"786B66F2",
x"7BDF68CB",
x"7F5D6A89",
x"82AB6C0C",
x"85A06D45",
x"882E6E33",
x"8A606EE4",
x"8C486F6C",
x"8E036FE4",
x"8FA9705F",
x"915370EE",
x"93077196",
x"94C67257",
x"96867329",
x"98357400",
x"99C274CE",
x"9B1B7588",
x"9C327626",
x"9D0476A2",
x"9D9576FF",
x"9DEE7741",
x"9E22776F",
x"9E427792",
x"9E6677B0",
x"9E9D77D2",
x"9EF377FE",
x"9F6E7834",
x"A00E7878",
x"A0C878CB",
x"A18E792C",
x"A2507998",
x"A2FA7A0B",
x"A3787A82",
x"A3BD7AF5",
x"A3C07B5B",
x"A37D7BAD",
x"A2F67BE1",
x"A2367BEF",
x"A14C7BD4",
x"A04A7B8F",
x"9F467B25",
x"9E547A9C",
x"9D8A7A02",
x"9CFA7968",
x"9CAE78E0",
x"9CAF7874",
x"9CFE7834",
x"9D957827",
x"9E69784E",
x"9F6778A3",
x"A07A791C",
x"A18879A9",
x"A2787A3A",
x"A3317ABC",
x"A39C7B20",
x"A3AE7B5A",
x"A3607B64",
x"A2B97B3D",
x"A1C67AED",
x"A0A57A7B",
x"9F7779F9",
x"9E637979",
x"9D92790F",
x"9D2878CA",
x"9D4078BD",
x"9DED78F4",
x"9F317977",
x"A1017A47",
x"A34C7B67",
x"A5F47CD0",
x"A8DC7E7A",
x"ABE48057",
x"AEF88261",
x"B20C8487",
x"B51686BF",
x"B81988F9",
x"BB198B2A",
x"BE1B8D43",
x"C11F8F39",
x"C41E9100",
x"C706928C",
x"C9C293D1",
x"CC3094C8",
x"CE34956C",
x"CFB495BE",
x"D09F95C2",
x"D0EE957F",
x"D0AF9504",
x"CFF5945F",
x"CEE293A3",
x"CD9B92DE",
x"CC439220",
x"CAF79173",
x"C9C790DF",
x"C8B99063",
x"C7C68FFA",
x"C6D68F9B",
x"C5D18F35",
x"C4998EBC",
x"C3138E1E",
x"C1338D52",
x"BEF08C4C",
x"BC568B10",
x"B97A89A1",
x"B67D8811",
x"B3878673",
x"B0C084DE",
x"AE4D8368",
x"AC458225",
x"AAAB8119",
x"A9738045",
x"A87B7F92",
x"A78F7EE8",
x"A66B7E1B",
x"A4CA7CFF",
x"A2647B6D",
x"9F047944",
x"9A8A7677",
x"94F3730B",
x"8E5D6F1C",
x"87076ADC",
x"7F4C668E",
x"7798627C",
x"705B5EE9",
x"6A035C14",
x"64EB5A28",
x"61515935",
x"5F525935",
x"5EE85A08",
x"5FEE5B7E",
x"62215D5C",
x"65335F60",
x"68C86156",
x"6C8D630E",
x"7035646D",
x"73896569",
x"76626606",
x"78AE6656",
x"7A6D6676",
x"7BAD6680",
x"7C816690",
x"7D0466BB",
x"7D50670D",
x"7D7A678A",
x"7D93682D",
x"7DA368EB",
x"7DB169B2",
x"7DBF6A72",
x"7DCB6B17",
x"7DD26B93",
x"7DD36BDC",
x"7DD06BEC",
x"7DCE6BC4",
x"7DCF6B68",
x"7DDC6AE5",
x"7DFD6A48",
x"7E3B69A0",
x"7E9768FA",
x"7F166865",
x"7FB267EB",
x"80676790",
x"812B6759",
x"81F46744",
x"82B8674C",
x"836F676F",
x"841367A8",
x"84A567F5",
x"852C6852",
x"85AE68C1",
x"86366942",
x"86D169D6",
x"87866A80",
x"88596B3B",
x"89496C04",
x"8A526CD5",
x"8B636DA3",
x"8C706E65",
x"8D656F12",
x"8E326FA3",
x"8ECD7014",
x"8F2E7068",
x"8F5670A1",
x"8F4D70CD",
x"8F2470F4",
x"8EE97121",
x"8EB1715F",
x"8E8D71B3",
x"8E8A721C",
x"8EAC7296",
x"8EF17317",
x"8F527392",
x"8FBB73F5",
x"901D7434",
x"90627440",
x"90797410",
x"905673A5",
x"8FF672FC",
x"8F5C7223",
x"8E957127",
x"8DB47019",
x"8CCD6F0D",
x"8BF76E19",
x"8B446D4D",
x"8AC16CB8",
x"8A736C63",
x"8A566C52",
x"8A606C7F",
x"8A816CDF",
x"8AA46D65",
x"8AB26DFD",
x"8A9F6E96",
x"8A606F1C",
x"89F06F80",
x"89556FBB",
x"889A6FCA",
x"87CF6FB0",
x"87066F76",
x"86506F29",
x"85BE6ED8",
x"85536E90",
x"85156E5B",
x"85006E3E",
x"85096E38",
x"85256E44",
x"85486E58",
x"85656E66",
x"85746E61",
x"85736E3D",
x"855D6DF0",
x"853A6D78",
x"85096CD5",
x"84D36C0C",
x"849E6B2A",
x"846D6A3A",
x"8442694E",
x"84206875",
x"840367BB",
x"83EC672E",
x"83D866D3",
x"83C466AD",
x"83AD66B7",
x"838A66E8",
x"83536731",
x"82FC677F",
x"827267BB",
x"81A167D1",
x"807967AB",
x"7EE5673A",
x"7CD96675",
x"7A556556",
x"775E63E9",
x"740A6238",
x"707C605D",
x"6CDC5E71",
x"69625C94",
x"663F5AE3",
x"63A7597A",
x"61C0586B",
x"60A657C5",
x"6064578C",
x"60F357BC",
x"6241584A",
x"642A5924",
x"66845A32",
x"69235B5F",
x"6BD85C95",
x"6E7A5DC1",
x"70EC5ED3",
x"73165FC2",
x"74EC6087",
x"766D6124",
x"779E619B",
x"788C61F4",
x"79446237",
x"79D36269",
x"7A4E6295",
x"7ABB62C2",
x"7B2562F4",
x"7B936331",
x"7C046377",
x"7C7963C8",
x"7CEA6423",
x"7D556483",
x"7DAF64E6",
x"7DF36545",
x"7E1A659E",
x"7E1E65E9",
x"7E016627",
x"7DC26652",
x"7D69666A",
x"7CFD6673",
x"7C8A666C",
x"7C1E6659",
x"7BC66641",
x"7B8E6627",
x"7B816610",
x"7BA16600",
x"7BEF65FA",
x"7C636601",
x"7CF66618",
x"7D98663E",
x"7E3C6672",
x"7ECF66B5",
x"7F486704",
x"7F9B675E",
x"7FC867BA",
x"7FCC6813",
x"7FB26862",
x"7F8068A1",
x"7F4468C9",
x"7F0668DB",
x"7ED268D4",
x"7EB068B8",
x"7EA06891",
x"7EA46866",
x"7EBA6845",
x"7EDB6834",
x"7F04683B",
x"7F31685C",
x"7F606891",
x"7F9368D4",
x"7FC96917",
x"8009694E",
x"8053696D",
x"80AE696F",
x"811A6951",
x"81946919",
x"821B68D5",
x"82A86896",
x"8332686C",
x"83B26866",
x"841E688D",
x"846D68E2",
x"849A695E",
x"849E69ED",
x"84796A7D",
x"842B6AF7",
x"83B96B48",
x"832A6B62",
x"82866B3F",
x"81D86AE8",
x"812B6A69",
x"808969DC",
x"7FFA6955",
x"7F8A68EC",
x"7F3868B2",
x"7F0A68AE",
x"7EFC68DF",
x"7F09693B",
x"7F2A69AD",
x"7F556A20",
x"7F816A80",
x"7FAA6ABB",
x"7FC56AC7",
x"7FD36AA1",
x"7FD66A51",
x"7FCF69E2",
x"7FC66965",
x"7FC268EB",
x"7FC86886",
x"7FDC683E",
x"7FFF681B",
x"802E681D",
x"8063683B",
x"8096686F",
x"80BC68AB",
x"80CF68E6",
x"80C76916",
x"80A06932",
x"80566938",
x"7FEA6923",
x"7F5968EF",
x"7EA0689A",
x"7DB56820",
x"7C93677F",
x"7B2866B1",
x"796C65B4",
x"77556487",
x"74E0632F",
x"721661B5",
x"6F066027",
x"6BCF5E94",
x"68995D11",
x"65925BB3",
x"62E95A8D",
x"60C859AC",
x"5F4F591B",
x"5E9258DA",
x"5E8D58E6",
x"5F345933",
x"606859B5",
x"61FD5A5A",
x"63C85B12",
x"659E5BCF",
x"67595C87",
x"68E15D31",
x"6A275DC8",
x"6B2B5E4C",
x"6BFA5EC1",
x"6CA35F24",
x"6D385F7C",
x"6DCF5FCB",
x"6E766013",
x"6F346059",
x"700D609E",
x"70FA60E6",
x"71F66135",
x"72F5618B",
x"73EA61EF",
x"74CF625C",
x"759B62D6",
x"764A6359",
x"76DB63E0",
x"774C6465",
x"77A164E2",
x"77D9654B",
x"77F9659B",
x"780065C9",
x"77F265CF",
x"77D265AA",
x"77A76559",
x"777664E2",
x"77486449",
x"7728639B",
x"772062E3",
x"77386235",
x"777961A1",
x"77E56139",
x"787F6110",
x"793F612E",
x"7A1D619B",
x"7B0C625A",
x"7BFD6363",
x"7CE064A7",
x"7DAA6610",
x"7E506786",
x"7ED268ED",
x"7F316A31",
x"7F796B3B",
x"7FBA6BFF",
x"80066C76",
x"80726CA7",
x"81106C9D",
x"81EC6C66",
x"830B6C19",
x"84676BC7",
x"85F46B83",
x"87986B58",
x"89396B4C",
x"8AB86B62",
x"8BF76B96",
x"8CDF6BE1",
x"8D656C38",
x"8D836C99",
x"8D436CF8",
x"8CBB6D54",
x"8C076DAA",
x"8B486DFA",
x"8A9D6E45",
x"8A226E8C",
x"89ED6ECE",
x"8A076F0A",
x"8A6D6F41",
x"8B136F70",
x"8BE06F93",
x"8CBB6FAB",
x"8D8A6FB7",
x"8E326FB7",
x"8EA46FB0",
x"8ED66FA1",
x"8ECB6F90",
x"8E8B6F7F",
x"8E286F70",
x"8DB56F66",
x"8D456F5F",
x"8CE96F5E",
x"8CAF6F5F",
x"8C9D6F65",
x"8CAF6F6E",
x"8CE56F79",
x"8D326F86",
x"8D8D6F94",
x"8DEA6FA1",
x"8E436FAB",
x"8E916FB0",
x"8ED06FAE",
x"8EFE6FA4",
x"8F1D6F92",
x"8F276F78",
x"8F1B6F58",
x"8EF66F35",
x"8EB16F16",
x"8E486EF9",
x"8DB66EE4",
x"8CFA6ED7",
x"8C176ED1",
x"8B136ECE",
x"89F36ECB",
x"88C56EBF",
x"87916EA4",
x"86606E72",
x"85356E21",
x"84106DAD",
x"82E96D0F",
x"81B76C45",
x"80696B51",
x"7EF66A34",
x"7D5268F3",
x"7B7A6799",
x"7973662E",
x"774B64C1",
x"7513635C",
x"72E8620E",
x"70E360E3",
x"6F205FE4",
x"6DB35F17",
x"6CAA5E81",
x"6C0D5E1F",
x"6BD85DF3",
x"6C025DF4",
x"6C7F5E21",
x"6D415E76",
x"6E3A5EED",
x"6F625F88",
x"70B56045",
x"72346124",
x"73DE6224",
x"75BA6346",
x"77C96487",
x"7A1165E5",
x"7C90675C",
x"7F4468E9",
x"82286A8D",
x"85386C45",
x"88726E16",
x"8BCB6FFE",
x"8F437202",
x"92D27421",
x"9670765A",
x"9A1078A3",
x"9DA57AF1",
x"A11C7D35",
x"A4637F59",
x"A767814F",
x"AA198302",
x"AC73846C",
x"AE6B8584",
x"B00F864C",
x"B16886CC",
x"B2878711",
x"B37E8729",
x"B45C8722",
x"B52C870A",
x"B5F486E6",
x"B6B386BC",
x"B761868B",
x"B7FA8653",
x"B8748612",
x"B8CF85C8",
x"B90C8578",
x"B939852E",
x"B96484F4",
x"B99F84D9",
x"B9FE84EA",
x"BA8C8535",
x"BB4E85BD",
x"BC3F8684",
x"BD4E877B",
x"BE658892",
x"BF6489AF",
x"C02F8AB8",
x"C0AB8B8D",
x"C0C78C1B",
x"C07F8C52",
x"BFDD8C2E",
x"BEF48BB8",
x"BDE78B05",
x"BCDD8A35",
x"BBFD896C",
x"BB6D88D0",
x"BB478887",
x"BB9E88A8",
x"BC6E8942",
x"BDAA8A50",
x"BF358BC3",
x"C0E48D79",
x"C2898F48",
x"C3F59101",
x"C4FF9276",
x"C5869382",
x"C57B9407",
x"C4D993FF",
x"C3B2936C",
x"C2209263",
x"C0519106",
x"BE728F7D",
x"BCB38DF1",
x"BB408C8B",
x"BA3C8B69",
x"B9B98A9B",
x"B9C08A29",
x"BA438A0D",
x"BB298A34",
x"BC4A8A84",
x"BD778AE0",
x"BE7F8B2C",
x"BF338B50",
x"BF6D8B39",
x"BF158AE2",
x"BE268A49",
x"BCAC897E",
x"BAC78894",
x"B8AB87A5",
x"B68E86CC",
x"B4B08625",
x"B34C85C3",
x"B28C85B5",
x"B28C85FD",
x"B34D8697",
x"B4BA8770",
x"B6A58871",
x"B8D4897E",
x"BB018A7A",
x"BCEA8B49",
x"BE568BD8",
x"BF208C18",
x"BF378C0A",
x"BEA28BB2",
x"BD788B1E",
x"BBDE8A5D",
x"B9FC8983",
x"B7F58898",
x"B5DA87A5",
x"B3AF86A2",
x"B15E8584",
x"AEC98436",
x"ABC2829F",
x"A81C80AB",
x"A3B87E46",
x"9E8A7B68",
x"98A2781F",
x"922E747E",
x"8B7470AB",
x"84D26CDB",
x"7EB16941",
x"79706614",
x"75666383",
x"72C961AD",
x"71B260A2",
x"72136064",
x"73BF60DD",
x"767061ED",
x"79D2636D",
x"7D906532",
x"815C6714",
x"84FD68F6",
x"88506AC4",
x"8B4F6C78",
x"8E016E13",
x"90816F9F",
x"92EF7126",
x"956472B4",
x"97F6744E",
x"9AA675F4",
x"9D6D779C",
x"A035793A",
x"A2DF7AC0",
x"A54D7C1E",
x"A7677D49",
x"A91C7E37",
x"AA6B7EEB",
x"AB5A7F68",
x"ABFA7FB9",
x"AC637FEA",
x"ACAB8008",
x"ACEA801F",
x"AD2E803C",
x"AD828066",
x"ADEA80A5",
x"AE6180FE",
x"AEE48174",
x"AF6E8208",
x"B00082BC",
x"B095838C",
x"B1338478",
x"B1E18576",
x"B2A1867B",
x"B377877D",
x"B466886C",
x"B56B893C",
x"B68289E2",
x"B7A38A53",
x"B8C78A90",
x"B9E78A98",
x"BAFE8A77",
x"BC088A38",
x"BD0789EA",
x"BDFE89A2",
x"BEF48970",
x"BFED8962",
x"C0ED8980",
x"C1F489D2",
x"C2FE8A58",
x"C4058B0D",
x"C4FE8BEC",
x"C5DA8CE9",
x"C68F8DFA",
x"C70F8F14",
x"C7589028",
x"C768912E",
x"C747921D",
x"C70292EA",
x"C6AD9390",
x"C65B9407",
x"C61E944C",
x"C606945F",
x"C61F943F",
x"C66793EF",
x"C6DA9378",
x"C76E92E2",
x"C8169241",
x"C8C991A2",
x"C979911A",
x"CA2590BC",
x"CAC99096",
x"CB6790B1",
x"CC049114",
x"CCA091B8",
x"CD3C9296",
x"CDCE939B",
x"CE4D94B3",
x"CEAA95C4",
x"CED896BA",
x"CECA9782",
x"CE7B980C",
x"CDEF9852",
x"CD359854",
x"CC649817",
x"CB9997AA",
x"CAF7971D",
x"CA9B9682",
x"CA9F95EF",
x"CB159576",
x"CC05952D",
x"CD6A951D",
x"CF31954F",
x"D14495C7",
x"D382967C",
x"D5C4975F",
x"D7E59859",
x"D9BA9951",
x"DB1F9A21",
x"DBF29AAE",
x"DC1F9ADC",
x"DB939A99",
x"DA5399DB",
x"D86798AB",
x"D5EA971D",
x"D2FC9548",
x"CFC69351",
x"CC689153",
x"C8FF8F67",
x"C5958D97",
x"C2208BDC",
x"BE858A22",
x"BA988846",
x"B6228623",
x"B0F08391",
x"AADA8074",
x"A3CD7CC1",
x"9BDA7883",
x"933273DB",
x"8A296EFF",
x"812B6A32",
x"78B565BE",
x"714161E9",
x"6B3E5EED",
x"66FD5CEE",
x"64AB5BFB",
x"644D5C08",
x"65BA5CF8",
x"68B05E9D",
x"6CD260BC",
x"71B76324",
x"76F965A0",
x"7C3B6809",
x"81346A44",
x"85AC6C42",
x"89886DFD",
x"8CBC6F78",
x"8F4D70B4",
x"914B71B7",
x"92C97289",
x"93DF7329",
x"94A4739D",
x"952973E5",
x"95847409",
x"95C2740C",
x"95EC73F9",
x"960E73DA",
x"962E73B7",
x"964D739A",
x"9670738B",
x"96947389",
x"96B87395",
x"96D573A7",
x"96EA73BD",
x"96F673CD",
x"96F673D5",
x"96EA73D4",
x"96D973CD",
x"96C273C3",
x"96AB73BE",
x"969873C7",
x"968B73E2",
x"968B7412",
x"969B7457",
x"96C274B0",
x"97087516",
x"97767586",
x"981375FC",
x"98E77678",
x"99F676F7",
x"9B3B777F",
x"9CAF7816",
x"9E4678C1",
x"9FEC7982",
x"A1887A5D",
x"A3077B4D",
x"A4567C4C",
x"A5677D4E",
x"A6387E49",
x"A6CA7F2D",
x"A7287FF4",
x"A7608091",
x"A77D8102",
x"A78E8147",
x"A7978161",
x"A7998159",
x"A7948135",
x"A77E8100",
x"A75480C2",
x"A7188081",
x"A6D28049",
x"A691801E",
x"A6708004",
x"A68A8001",
x"A6FD8016",
x"A7DD8047",
x"A9368092",
x"AB0280F7",
x"AD28816E",
x"AF8781F4",
x"B1EB8280",
x"B4218307",
x"B5F88382",
x"B74D83EC",
x"B80A843D",
x"B82F8476",
x"B7CF8495",
x"B708849E",
x"B6048495",
x"B4EB847D",
x"B3DD8459",
x"B2EE8429",
x"B22383ED",
x"B16E839F",
x"B0B8833C",
x"AFE682C0",
x"AEDC8226",
x"AD898171",
x"ABF080A5",
x"AA1E7FC7",
x"A8357EEB",
x"A6637E1C",
x"A4DE7D6F",
x"A3D67CFA",
x"A3737CCA",
x"A3C77CEF",
x"A4D07D6B",
x"A6747E3D",
x"A8847F54",
x"AAC3809F",
x"ACEE8200",
x"AEC48356",
x"B0168481",
x"B0C28562",
x"B0BD85E3",
x"B01685F4",
x"AEE78594",
x"AD5984C5",
x"AB958398",
x"A9BD821F",
x"A7E38070",
x"A60B7E9C",
x"A4217CB0",
x"A2077AB2",
x"9F9278A0",
x"9C9B7678",
x"99057431",
x"94C871C8",
x"8FF06F43",
x"8AAA6CAA",
x"85386A16",
x"7FF067A4",
x"7B2F657A",
x"775163BE",
x"749E6291",
x"734B620D",
x"736D623C",
x"74FA631D",
x"77CB649D",
x"7B9D669B",
x"802568F5",
x"850D6B7D",
x"8A076E0A",
x"8ECD7078",
x"932C72AD",
x"97017496",
x"9A3B762C",
x"9CD2776E",
x"9ED07862",
x"A03E7912",
x"A1297988",
x"A19F79CA",
x"A1AB79E1",
x"A15679D6",
x"A0AE79A9",
x"9FBC7962",
x"9E8F7908",
x"9D39789D",
x"9BCC782D",
x"9A5D77BE",
x"99007758",
x"97C67703",
x"96C176C4",
x"95F6769F",
x"956E7695",
x"952C76A5",
x"952B76CA",
x"95667702",
x"95D37747",
x"96697790",
x"971877DA",
x"97D2781C",
x"98877853",
x"99247875",
x"9998787F",
x"99D6786B",
x"99D37833",
x"998877D7",
x"98F67754",
x"982576AA",
x"971F75E1",
x"95FC74FE",
x"94CC740D",
x"93AA7320",
x"92AA7248",
x"91DC7195",
x"914C7119",
x"910170DF",
x"90FB70EF",
x"91327148",
x"919D71E1",
x"922972A7",
x"92C97386",
x"936A7464",
x"93FB7529",
x"946D75BE",
x"94B57615",
x"94C87629",
x"94A175F9",
x"943F7593",
x"93A77503",
x"92E2745C",
x"91FB73AF",
x"91047309",
x"90117274",
x"8F3271F0",
x"8E7A7180",
x"8DFA7120",
x"8DBB70CB",
x"8DC67080",
x"8E1A7044",
x"8EB2701C",
x"8F867010",
x"9087702D",
x"91A5707C",
x"92D07102",
x"93F971BD",
x"950D72A1",
x"960073A1",
x"96C674A5",
x"97567592",
x"97A97650",
x"97BB76CD",
x"978A76FE",
x"971876DE",
x"966D767B",
x"959475E2",
x"949E752F",
x"93A47479",
x"92C073E1",
x"92137379",
x"91BC7355",
x"91D9737B",
x"927E73EA",
x"93B6749C",
x"957D7581",
x"97BC7689",
x"9A5277A0",
x"9D0B78B3",
x"9FAF79B2",
x"A2037A8E",
x"A3D07B3C",
x"A4F17BB7",
x"A5537BFC",
x"A4F77C0E",
x"A3F67BEE",
x"A2777BA3",
x"A0B27B36",
x"9EDC7AAC",
x"9D227A0C",
x"9BA1795A",
x"9A5F7895",
x"994977B6",
x"983976B4",
x"96F37582",
x"9539740F",
x"92D0724E",
x"8F8A7034",
x"8B566DBE",
x"863F6AF6",
x"806F67ED",
x"7A2D64C5",
x"73D261A1",
x"6DC45EB1",
x"68605C1E",
x"63FF5A11",
x"60DA58A6",
x"5F0D57EE",
x"5E9E57E7",
x"5F6E5884",
x"614A59AB",
x"63EF5B38",
x"67165D08",
x"6A765EF7",
x"6DD460E7",
x"70FC62C1",
x"73D26474",
x"764665FC",
x"78586755",
x"7A136883",
x"7B8D6987",
x"7CDC6A69",
x"7E1B6B2A",
x"7F606BCF",
x"80BE6C5E",
x"82426CD9",
x"83F36D4E",
x"85CF6DC1",
x"87CF6E3E",
x"89E66ECE",
x"8C016F73",
x"8E0B702D",
x"8FF070F2",
x"919871B4",
x"92F77264",
x"940072EB",
x"94B17339",
x"95087341",
x"95107300",
x"94D2727E",
x"945771C7",
x"93B170F5",
x"92E37020",
x"91F96F61",
x"90F46ECB",
x"8FDC6E6E",
x"8EB16E48",
x"8D7B6E54",
x"8C456E85",
x"8B1A6EC5",
x"8A096F05",
x"89256F34",
x"88806F4D",
x"88276F4A",
x"88246F37",
x"88776F1C",
x"891B6F09",
x"8A046F0A",
x"8B1E6F27",
x"8C556F62",
x"8D916FB7",
x"8EBC701C",
x"8FC57082",
x"909F70DE",
x"91427124",
x"91AB7154",
x"91DA716B",
x"91D67174",
x"91A47176",
x"914C7180",
x"90D8719D",
x"905271D4",
x"8FC57224",
x"8F3C728A",
x"8EC172F8",
x"8E597362",
x"8E0A73B6",
x"8DD373E5",
x"8DAE73E5",
x"8D9273B0",
x"8D737344",
x"8D4372A6",
x"8CF371DC",
x"8C7D70F6",
x"8BDA6FFC",
x"8B0E6EFE",
x"8A276E05",
x"89316D1D",
x"88426C51",
x"876D6BA7",
x"86C56B26",
x"86526AD1",
x"86176AA7",
x"860B6AA6",
x"86226AC7",
x"86436AFD",
x"865B6B3B",
x"864F6B6F",
x"86146B89",
x"85A06B79",
x"84F66B35",
x"84216ABD",
x"83356A10",
x"8248693C",
x"81726852",
x"80C36765",
x"804B668D",
x"800D65DF",
x"80036566",
x"8020652F",
x"804E6537",
x"80796577",
x"808C65E2",
x"80706662",
x"801D66E2",
x"7F8A674C",
x"7EBB6791",
x"7DB567A4",
x"7C86677D",
x"7B37671B",
x"79D56683",
x"786765BE",
x"76F064D6",
x"756F63D6",
x"73DE62C9",
x"723461B8",
x"706960A9",
x"6E795FA4",
x"6C625EA8",
x"6A2A5DBB",
x"67DF5CDD",
x"65975C14",
x"636F5B61",
x"61875ACD",
x"5FFF5A5A",
x"5EF35A0E",
x"5E7C59EE",
x"5EA359FB",
x"5F6B5A36",
x"60C55A9B",
x"629D5B22",
x"64D15BC2",
x"673E5C71",
x"69BC5D21",
x"6C2E5DCB",
x"6E795E63",
x"708C5EE7",
x"72635F5A",
x"74075FC3",
x"7584602B",
x"76F0609E",
x"7860612D",
x"79E861E0",
x"7B9062BF",
x"7D5C63CB",
x"7F4864FC",
x"81416645",
x"832F6796",
x"84FB68D8",
x"868A69F9",
x"87C36AEB",
x"889E6BA3",
x"89136C21",
x"892B6C6F",
x"88F76C99",
x"88906CB1",
x"88146CCB",
x"87A16CF9",
x"87516D47",
x"87356DB7",
x"87556E47",
x"87AC6EE9",
x"882B6F8A",
x"88B87017",
x"89357079",
x"8981709F",
x"8981707C",
x"8922700F",
x"885C6F5E",
x"87386E79",
x"85C86D75",
x"842E6C6C",
x"82916B7C",
x"811A6ABA",
x"7FF26A38",
x"7F346A04",
x"7EF16A1D",
x"7F2E6A7D",
x"7FDC6B11",
x"80DF6BC8",
x"82156C86",
x"83586D33",
x"847D6DBA",
x"85656E0C",
x"85F96E20",
x"862E6DF6",
x"86046D94",
x"858A6D09",
x"84D56C66",
x"83FC6BBE",
x"831B6B24",
x"824E6AA8",
x"81A86A58",
x"813C6A38",
x"81136A4E",
x"81316A97",
x"81986B0F",
x"82436BAB",
x"832B6C63",
x"84486D2E",
x"858A6DFF",
x"86E66ECE",
x"884C6F93",
x"89A87047",
x"8AED70E4",
x"8C067168",
x"8CE571CF",
x"8D80721A",
x"8DCF7243",
x"8DD2724A",
x"8D8B722B",
x"8D0871E6",
x"8C56717B",
x"8B8470EB",
x"8AA4703A",
x"89C36F72",
x"88F06E9E",
x"88326DD1",
x"878B6D19",
x"86FD6C87",
x"86866C2B",
x"86206C0C",
x"85C96C2A",
x"857D6C7D",
x"85386CF6",
x"84FB6D80",
x"84C46E00",
x"84906E5C",
x"845C6E80",
x"84246E5B",
x"83DD6DE8",
x"83836D2D",
x"830A6C38",
x"826D6B20",
x"81AA69FD",
x"80C268E8",
x"7FBE67F7",
x"7EA8673B",
x"7D9366B7",
x"7C8B6669",
x"7BA36648",
x"7ADF6641",
x"7A41663E",
x"79C2662B",
x"795365F3",
x"78DC6587",
x"784264E0",
x"776F63FF",
x"764C62E6",
x"74CF61A7",
x"72FC6053",
x"70DE5F01",
x"6E905DC6",
x"6C375CBB",
x"69FC5BEE",
x"68095B6E",
x"66865B3F",
x"65905B5D",
x"653B5BC2",
x"658D5C5D",
x"66805D1C",
x"68005DEE",
x"69F65EC3",
x"6C425F90",
x"6EC7604F",
x"71686104",
x"740C61B7",
x"76A56273",
x"792A6349",
x"7B936442",
x"7DE56569",
x"802066BE",
x"8249683B",
x"846669D2",
x"867A6B72",
x"88846D03",
x"8A7E6E6E",
x"8C656FA0",
x"8E2A7089",
x"8FC67120",
x"912E7165",
x"9258715F",
x"9342711D",
x"93F070B1",
x"946A7031",
x"94C16FB5",
x"95076F4F",
x"95566F12",
x"95BE6F05",
x"964B6F29",
x"96FB6F7A",
x"97BF6FE9",
x"98777064",
x"98F770CE",
x"990E7112",
x"98877113",
x"973570C1",
x"94FE700F",
x"91DF6EFC",
x"8DEC6D8F",
x"89526BDE",
x"845669FF",
x"7F486814",
x"7A7C663C",
x"763C6494",
x"72C76332",
x"703E6224",
x"6EAD6170",
x"6E076113",
x"6E2D6101",
x"6EED612B",
x"70196181",
x"717A61F0",
x"72E9626A",
x"744562E4",
x"75776356",
x"767563BE",
x"7737641B",
x"77C2646F",
x"781864BC",
x"783F6509",
x"783E6555",
x"781A65A4",
x"77DB65F5",
x"77866645",
x"77236690",
x"76B266CE",
x"763466F5",
x"75A466F9",
x"74F966CF",
x"742A6670",
x"733465D9",
x"7218650D",
x"70E16418",
x"6FA7630D",
x"6E936207",
x"6DD46128",
x"6DA16090",
x"6E30605D",
x"6FA760A8",
x"721D6179",
x"758D62D0",
x"79D8649B",
x"7EC266BF",
x"83FD6914",
x"892E6B70",
x"8DF76DA7",
x"92096F96",
x"95257120",
x"972B7237",
x"981472DA",
x"97FB7313",
x"971172F9",
x"959572A4",
x"93CD7234",
x"91FD71C0",
x"905C715E",
x"8F117117",
x"8E2E70F0",
x"8DB470E5",
x"8D9070E8",
x"8DA770EB",
x"8DD770DE",
x"8E0170B5",
x"8E0B706C",
x"8DE97000",
x"8D926F78",
x"8D126EDF",
x"8C796E47",
x"8BD86DBB",
x"8B406D4A",
x"8ABE6CF8",
x"8A506CC5",
x"89EC6CA8",
x"89776C92",
x"88CE6C69",
x"87C66C16",
x"863B6B82",
x"84096A94",
x"811A6944",
x"7D6D678C",
x"79176573",
x"7439630D",
x"6F0F6074",
x"69D85DC9",
x"64DF5B33",
x"606858D7",
x"5CB056D4",
x"59DF5546",
x"5813543F",
x"574D53C3",
x"577E53CE",
x"58885451",
x"5A3E5535",
x"5C72565A",
x"5EF057A1",
x"618A58E6",
x"64175A10",
x"66795B04",
x"689A5BB8",
x"6A725C25",
x"6BFD5C56",
x"6D445C57",
x"6E4F5C3F",
x"6F315C2B",
x"6FF75C31",
x"70B25C69",
x"716F5CE3",
x"72345DA7",
x"73065EAE",
x"73E25FED",
x"74BF614E",
x"759162B5",
x"76466403",
x"76D1651B",
x"772165E5",
x"772B664E",
x"76EC664F",
x"766565E8",
x"75A36525",
x"74B56417",
x"73B162D6",
x"72AD617D",
x"71BC6025",
x"70F05EE3",
x"70545DC9",
x"6FEC5CE4",
x"6FB45C36",
x"6FA85BC2",
x"6FBE5B81",
x"6FEB5B6B",
x"70275B7A",
x"706F5BA5",
x"70BE5BE9",
x"711A5C40",
x"71845CAE",
x"72025D31",
x"72935DCB",
x"73385E7C",
x"73EA5F3F",
x"74A06011",
x"754B60EC",
x"75DC61C3",
x"7645628B",
x"767C633B",
x"767D63C8",
x"7646642A",
x"75E3645C",
x"75606460",
x"74CF643B",
x"744463EF",
x"73D26389",
x"738A6311",
x"73796295",
x"73A0621F",
x"740061BB",
x"7491616F",
x"75486145",
x"76146142",
x"76E66164",
x"77AD61AD",
x"78596213",
x"78DF628D",
x"7935630E",
x"7958638B",
x"794263F3",
x"78F96439",
x"78806458",
x"77E0644B",
x"77276414",
x"766563BE",
x"75AB6356",
x"750C62EF",
x"749A629B",
x"7463626D",
x"74736273",
x"74CE62B5",
x"75726335",
x"765563F0",
x"776B64DA",
x"78A065E3",
x"79DD66FA",
x"7B10680D",
x"7C256909",
x"7D1169E1",
x"7DCC6A8A",
x"7E536AFF",
x"7EAB6B3B",
x"7ED96B45",
x"7EE66B1D",
x"7ED96ACC",
x"7EBB6A5C",
x"7E9069D2",
x"7E59693C",
x"7E1668A6",
x"7DC86814",
x"7D6F6794",
x"7D09672D",
x"7C9966E0",
x"7C2066B1",
x"7B9E669A",
x"7B136694",
x"7A796690",
x"79C96680",
x"78FA6652",
x"77FD65F6",
x"76C56562",
x"7547648A",
x"737D6373",
x"716C6221",
x"6F1E60A7",
x"6CAE5F1A",
x"6A3A5D91",
x"67EB5C2B",
x"65EB5AFE",
x"64635A1F",
x"6378599B",
x"633D5977",
x"63BD59AF",
x"64F05A3B",
x"66C45B07",
x"69135C01",
x"6BB25D17",
x"6E765E32",
x"712E5F45",
x"73B46042",
x"75E96127",
x"77BC61ED",
x"79286298",
x"7A32632F",
x"7AEC63B5",
x"7B696431",
x"7BC264AA",
x"7C0E6523",
x"7C62659E",
x"7CC9661D",
x"7D4C66A0",
x"7DED6727",
x"7EA867AE",
x"7F766837",
x"804968BF",
x"811B6945",
x"81DF69C9",
x"828D6A47",
x"831D6ABA",
x"838A6B1E",
x"83D26B6F",
x"83F46BA1",
x"83F06BAE",
x"83C86B93",
x"837F6B49",
x"83186AD7",
x"829A6A3F",
x"82096990",
x"816D68D8",
x"80CE682B",
x"80356799",
x"7FAB6731",
x"7F3A66FC",
x"7EE766FD",
x"7EBF6732",
x"7EC56793",
x"7EFC6811",
x"7F6368A0",
x"7FFA6934",
x"80BC69C4",
x"81A16A4E",
x"82A36AD2",
x"83B56B58",
x"84D26BE3",
x"85EF6C7A",
x"87066D1E",
x"880E6DCD",
x"89046E78",
x"89E26F14",
x"8AA26F90",
x"8B426FDB",
x"8BBE6FE6",
x"8C136FAB",
x"8C3C6F2E",
x"8C3C6E75",
x"8C116D92",
x"8BBE6C99",
x"8B456BA0",
x"8AAB6ABD",
x"89FA69FD",
x"8938696D",
x"88706910",
x"87AB68E5",
x"86F768E5",
x"865F6907",
x"85ED6948",
x"85AB699E",
x"85A26A04",
x"85D36A79",
x"863F6AF9",
x"86E06B83",
x"87AB6C13",
x"88906CA3",
x"89796D2B",
x"8A526DA3",
x"8B046E00",
x"8B806E3A",
x"8BB96E4D",
x"8BAF6E33",
x"8B676DF3",
x"8AF36D93",
x"8A676D1D",
x"89E06CA3",
x"89796C30",
x"89456BD5",
x"89566B9E",
x"89B26B96",
x"8A556BC1",
x"8B316C20",
x"8C316CB3",
x"8D3F6D70",
x"8E426E52",
x"8F256F4A",
x"8FD8704A",
x"904D7141",
x"9083721F",
x"907672D1",
x"902C734A",
x"8FA97379",
x"8EF4735A",
x"8E1472E5",
x"8D0D7220",
x"8BE67114",
x"8AA16FD1",
x"89426E69",
x"87CB6CF0",
x"86366B7A",
x"84836A14",
x"82A768C5",
x"8093678C",
x"7E3A6660",
x"7B8D6532",
x"788463F3",
x"75206291",
x"716C6104",
x"6D845F49",
x"69965D6A",
x"65D55B81",
x"628059A8",
x"5FD85805",
x"5E0F56BC",
x"5D4D55EB",
x"5D9D55A8",
x"5EF855F4",
x"613A56CA",
x"642D5811",
x"678C59A5",
x"6B115B60",
x"6E7A5D18",
x"71945EAC",
x"743E6006",
x"766D6117",
x"782D61E4",
x"7991627D",
x"7AB962F7",
x"7BC6636C",
x"7CD563F2",
x"7DF5649E",
x"7F2C657A",
x"80796687",
x"81D267BC",
x"8328690D",
x"84736A65",
x"85AA6BB1",
x"86CF6CE2",
x"87EA6DE9",
x"89076EBE",
x"8A316F5F",
x"8B766FCF",
x"8CDA7016",
x"8E62703A",
x"90047048",
x"91BB704D",
x"93747054",
x"95257069",
x"96C17099",
x"983B70EB",
x"998F7165",
x"9ABE720C",
x"9BC272DB",
x"9CA273CE",
x"9D5F74DA",
x"9DFB75EB",
x"9E7876F4",
x"9EDC77E0",
x"9F2B789F",
x"9F6D7926",
x"9FAF796F",
x"A0007982",
x"A06E7968",
x"A10A7934",
x"A1DC78FC",
x"A2E778D7",
x"A42678D6",
x"A58A7908",
x"A6FB796F",
x"A85F7A06",
x"A9957AC3",
x"AA857B8E",
x"AB1F7C51",
x"AB597CFA",
x"AB397D74",
x"AAD37DB7",
x"AA3D7DC1",
x"A99B7D99",
x"A9077D4A",
x"A89E7CE4",
x"A86E7C7B",
x"A87E7C1B",
x"A8C37BD1",
x"A92E7BA0",
x"A9A17B89",
x"AA027B84",
x"AA367B88",
x"AA297B89",
x"A9CD7B7F",
x"A9217B60",
x"A82B7B29",
x"A6F87AD7",
x"A59C7A6E",
x"A42679EE",
x"A2A6795D",
x"A12978C0",
x"9FB6781B",
x"9E537772",
x"9D0076C8",
x"9BC07625",
x"9A95758D",
x"99847506",
x"98957499",
x"97CF744B",
x"97367421",
x"96D0741A",
x"969D7433",
x"96957462",
x"96AE749D",
x"96D974D4",
x"970174F5",
x"971A74F5",
x"971474CA",
x"96E47472",
x"968A73F2",
x"96067351",
x"955F72A1",
x"949C71F0",
x"93C87151",
x"92EA70CD",
x"920A706B",
x"9129702D",
x"904B700C",
x"8F736FFC",
x"8EA46FF0",
x"8DE06FDC",
x"8D316FB4",
x"8C9A6F6E",
x"8C206F06",
x"8BBE6E7D",
x"8B6F6DD7",
x"8B216D16",
x"8ABC6C3E",
x"8A246B52",
x"89356A54",
x"87D5693E",
x"85EC6813",
x"837266D2",
x"8070657F",
x"7D016420",
x"794E62C1",
x"758D6170",
x"71FF6041",
x"6EDF5F41",
x"6C685E83",
x"6AC25E12",
x"6A075DF4",
x"6A3E5E2C",
x"6B5B5EB3",
x"6D445F86",
x"6FD26098",
x"72DE61E2",
x"763E635C",
x"79CF6503",
x"7D7766D2",
x"812568CB",
x"84D36AEC",
x"88806D31",
x"8C2E6F94",
x"8FDF720A",
x"93927482",
x"974276E8",
x"9AE17925",
x"9E5A7B23",
x"A1977CCE",
x"A47A7E19",
x"A6EA7EFE",
x"A8D07F78",
x"AA1E7F98",
x"AACA7F67",
x"AADA7EFB",
x"AA577E68",
x"A9567DC0",
x"A7F17D15",
x"A6497C71",
x"A4807BDD",
x"A2B97B5D",
x"A11A7AF4",
x"9FC37AA3",
x"9ED37A6F",
x"9E667A61",
x"9E8F7A81",
x"9F597ADB",
x"A0C87B7C",
x"A2D37C6F",
x"A5677DB7",
x"A8697F4F",
x"ABAF812F",
x"AF0E8343",
x"B25C8570",
x"B56A8797",
x"B816899A",
x"BA478B5C",
x"BBF18CC8",
x"BD168DCF",
x"BDC98E70",
x"BE258EAF",
x"BE498E9D",
x"BE5B8E4B",
x"BE7B8DD3",
x"BEC08D4C",
x"BF398CC9",
x"BFE68C5D",
x"C0BD8C11",
x"C1AC8BE7",
x"C29B8BDD",
x"C36E8BED",
x"C4158C0A",
x"C47E8C25",
x"C4A38C36",
x"C48C8C32",
x"C4448C14",
x"C3DE8BD9",
x"C3718B88",
x"C3128B2B",
x"C2D08ACC",
x"C2B98A7B",
x"C2CD8A46",
x"C3058A35",
x"C3548A4C",
x"C3A88A85",
x"C3E88AD8",
x"C4018B32",
x"C3E48B80",
x"C3898BAE",
x"C2F28BAC",
x"C22A8B73",
x"C1438AFE",
x"C0548A59",
x"BF788992",
x"BEC688C2",
x"BE4F87FE",
x"BE19875D",
x"BE2886F3",
x"BE6B86C6",
x"BED486D9",
x"BF4A8722",
x"BFB78797",
x"C0098824",
x"C03688B8",
x"C03A8946",
x"C01C89C3",
x"BFE48A29",
x"BFA38A77",
x"BF648AAE",
x"BF2B8ACC",
x"BEF48AD2",
x"BEB08ABE",
x"BE4D8A8A",
x"BDAA8A2E",
x"BCB289A4",
x"BB4E88E7",
x"B97587F9",
x"B72D86DC",
x"B48C859B",
x"B1B58445",
x"AECF82E7",
x"AC088192",
x"A97E804D",
x"A7457F19",
x"A55C7DF4",
x"A3A87CC7",
x"A1FD7B81",
x"A01C7A03",
x"9DC57839",
x"9AB9760B",
x"96CD736C",
x"91ED7062",
x"8C276CF9",
x"85A5694E",
x"7EB26586",
x"77AE61CE",
x"71005E56",
x"6B0D5B4C",
x"662B58D0",
x"629656FF",
x"606C55E3",
x"5FA75578",
x"602455B2",
x"61A95675",
x"63EB57A4",
x"669B591A",
x"69735AB6",
x"6C345C5C",
x"6EB75DF0",
x"70E65F60",
x"72BD60A4",
x"744761B4",
x"75996293",
x"76C96344",
x"77F263CF",
x"791E6441",
x"7A5964A0",
x"7BA364F6",
x"7CF2654C",
x"7E3B65AA",
x"7F706611",
x"80836687",
x"8168670A",
x"82156796",
x"828A6826",
x"82C268B2",
x"82C46937",
x"829769AB",
x"82456A0D",
x"81DB6A58",
x"81656A8C",
x"80F46AA8",
x"80946AB4",
x"80526AB0",
x"80356AA0",
x"80446A8C",
x"807E6A75",
x"80E06A62",
x"81636A54",
x"81FA6A51",
x"82986A5C",
x"83346A7A",
x"83C26AB0",
x"843C6AFC",
x"84A26B62",
x"84F96BDE",
x"85486C6B",
x"859B6CFD",
x"85FE6D8A",
x"867D6E08",
x"871A6E65",
x"87D96E9C",
x"88B16EA7",
x"89976E86",
x"8A796E3D",
x"8B456DD8",
x"8BE76D63",
x"8C556CEE",
x"8C846C86",
x"8C776C37",
x"8C396C07",
x"8BD96BFC",
x"8B6F6C13",
x"8B136C48",
x"8AD96C99",
x"8AD66CFA",
x"8B106D6C",
x"8B876DE5",
x"8C2F6E63",
x"8CFA6EDE",
x"8DCC6F51",
x"8E8E6FB1",
x"8F286FF8",
x"8F887017",
x"8FA27009",
x"8F776FC4",
x"8F0B6F47",
x"8E6F6E96",
x"8DAF6DBB",
x"8CE36CCA",
x"8C1D6BD7",
x"8B676AF7",
x"8ACF6A45",
x"8A5569D2",
x"89F969A7",
x"89B569C8",
x"89816A2D",
x"89586AC9",
x"89326B89",
x"890E6C54",
x"88EF6D14",
x"88D56DB5",
x"88C86E2B",
x"88C96E6E",
x"88DF6E7D",
x"89086E62",
x"89466E27",
x"89936DDC",
x"89EA6D90",
x"8A486D4F",
x"8AA46D24",
x"8AFD6D14",
x"8B4F6D20",
x"8B986D42",
x"8BD96D73",
x"8C116DAB",
x"8C3F6DDF",
x"8C636E08",
x"8C796E20",
x"8C7B6E29",
x"8C666E21",
x"8C2F6E10",
x"8BCE6DF9",
x"8B366DDF",
x"8A5D6DBF",
x"89356D96",
x"87B26D58",
x"85C56CF8",
x"83656C65",
x"808E6B90",
x"7D426A6B",
x"798E68F0",
x"75876721",
x"714E650B",
x"6D0D62C2",
x"68F6605F",
x"653B5E03",
x"620D5BC9",
x"5F9259D2",
x"5DE5582F",
x"5D1456F3",
x"5D1C5622",
x"5DE855BF",
x"5F5B55C4",
x"614E5626",
x"639656DD",
x"660D57D9",
x"6890590F",
x"6B065A74",
x"6D5C5BFA",
x"6F8C5D94",
x"71915F35",
x"737060CC",
x"752D624E",
x"76CB63AE",
x"784E64E2",
x"79B865E5",
x"7B0D66B8",
x"7C4E675F",
x"7D7C67E5",
x"7E9A6855",
x"7FAE68BB",
x"80BC6923",
x"81CB6994",
x"82DC6A14",
x"83F36AA0",
x"850D6B34",
x"86256BCA",
x"87356C59",
x"88326CDC",
x"89146D52",
x"89D06DB7",
x"8A5F6E12",
x"8ABC6E62",
x"8AE96EB1",
x"8AE76F02",
x"8ABF6F52",
x"8A7C6FA3",
x"8A2C6FEE",
x"89DD702B",
x"89A27054",
x"898A705F",
x"899F704B",
x"89EF701A",
x"8A7A6FD2",
x"8B456F82",
x"8C4B6F3A",
x"8D836F0A",
x"8EE26F08",
x"905C6F3E",
x"91E36FB4",
x"936C706C",
x"94EA715C",
x"96597275",
x"97AE73A1",
x"98E774CA",
x"99FE75D4",
x"9AF376AD",
x"9BC27744",
x"9C6A7790",
x"9CEC7795",
x"9D487757",
x"9D8076E8",
x"9D9C765E",
x"9DA275CB",
x"9D9B7548",
x"9D9074E5",
x"9D8274B0",
x"9D7874AA",
x"9D6E74D2",
x"9D60751F",
x"9D45757E",
x"9D1475DC",
x"9CC3762A",
x"9C4F7654",
x"9BB8764E",
x"9B077615",
x"9A4975AA",
x"99917515",
x"98F77467",
x"988F73AD",
x"986972FE",
x"988B7268",
x"98F671FB",
x"999A71BA",
x"9A6371A7",
x"9B3471BE",
x"9BEC71F2",
x"9C6D7234",
x"9C9A7272",
x"9C63729F",
x"9BC072AB",
x"9AB67290",
x"9955724B",
x"97B571DF",
x"95F7715A",
x"943C70C4",
x"92AA7034",
x"915A6FB7",
x"90646F5F",
x"8FD66F33",
x"8FAF6F38",
x"8FE46F6B",
x"90626FC1",
x"910E702A",
x"91CA7094",
x"927A70E9",
x"9303711C",
x"9355711D",
x"936570EB",
x"93347088",
x"92C96FFE",
x"922C6F5B",
x"916C6EB0",
x"908B6E08",
x"8F8D6D6E",
x"8E696CE1",
x"8D106C58",
x"8B6F6BCA",
x"89706B20",
x"87066A49",
x"84286937",
x"80E067E3",
x"7D486652",
x"79846494",
x"75CE62C2",
x"725B6101",
x"6F6B5F73",
x"6D2D5E3C",
x"6BCB5D77",
x"6B575D33",
x"6BCF5D76",
x"6D215E33",
x"6F2A5F55",
x"71BA60BC",
x"74A06249",
x"77AD63DC",
x"7AB86559",
x"7DA166AD",
x"805567CF",
x"82CC68BE",
x"85096984",
x"87116A2D",
x"88ED6AC9",
x"8AA86B69",
x"8C496C1A",
x"8DD26CE2",
x"8F436DC5",
x"909D6EC1",
x"91D86FCE",
x"92F070DE",
x"93E571E6",
x"94B572D8",
x"956273AA",
x"95F37451",
x"966D74CB",
x"96DC751A",
x"974B7546",
x"97C37558",
x"98507561",
x"98FA756C",
x"99C5758C",
x"9AB575C8",
x"9BC97627",
x"9CFD76AA",
x"9E49774A",
x"9FA977FE",
x"A11478B9",
x"A2857971",
x"A3FA7A1C",
x"A5717AB3",
x"A6EE7B36",
x"A8777BA9",
x"AA0E7C13",
x"ABB67C81",
x"AD717CFA",
x"AF397D84",
x"B1047E25",
x"B2C57EDA",
x"B4687F99",
x"B5E0805E",
x"B7188118",
x"B80781BC",
x"B8A68240",
x"B8FB829E",
x"B90B82D4",
x"B8E882E6",
x"B8A582DA",
x"B85682BD",
x"B80C829B",
x"B7DA827E",
x"B7C98271",
x"B7DD827E",
x"B81982A9",
x"B87B82F4",
x"B8FE8361",
x"B99E83ED",
x"BA578497",
x"BB268557",
x"BC0C862B",
x"BD05870B",
x"BE1487F1",
x"BF3288D6",
x"C05D89B2",
x"C18E8A7D",
x"C2B78B2F",
x"C3D18BC5",
x"C4CA8C38",
x"C5988C86",
x"C62A8CAF",
x"C6788CB5",
x"C67A8C9D",
x"C6298C69",
x"C58B8C20",
x"C4A08BC8",
x"C3748B67",
x"C2118B00",
x"C0878A94",
x"BEE48A25",
x"BD3A89B2",
x"BB988939",
x"BA0988B9",
x"B89B8835",
x"B75187AC",
x"B6368727",
x"B54E86A8",
x"B49C863C",
x"B42385E9",
x"B3E785B6",
x"B3E385A9",
x"B41185BD",
x"B46885EC",
x"B4D68627",
x"B543865A",
x"B5968674",
x"B5B5865E",
x"B5888611",
x"B5028584",
x"B42284BF",
x"B2F483D6",
x"B19282E1",
x"B0228201",
x"AECC8154",
x"ADB380F0",
x"ACF080DB",
x"AC7D810F",
x"AC45816E",
x"AC1481CA",
x"ABA281EB",
x"AA9B8194",
x"A8AC808B",
x"A5957EAD",
x"A1327BE5",
x"9B837840",
x"94B573DF",
x"8D1E6F08",
x"85346A04",
x"7D7A6531",
x"767960E2",
x"70A85D5F",
x"6C5F5ADD",
x"69CE5975",
x"68F75928",
x"69B759DD",
x"6BC55B66",
x"6EC85D8B",
x"725D600E",
x"762E62B7",
x"79ED6552",
x"7D6A67B8",
x"808C69D4",
x"834F6B99",
x"85C26D0A",
x"87FD6E31",
x"8A176F1D",
x"8C276FE1",
x"8E35708D",
x"90467131",
x"924F71D5",
x"94457282",
x"96157337",
x"97B273F5",
x"991474B9",
x"9A38757E",
x"9B22763E",
x"9BE376FC",
x"9C8777B2",
x"9D247861",
x"9DC8790C",
x"9E8179B4",
x"9F597A5D",
x"A04D7B04",
x"A15D7BAC",
x"A27D7C51",
x"A3A27CF2",
x"A4C07D89",
x"A5CA7E14",
x"A6B67E8E",
x"A77F7EF5",
x"A8227F47",
x"A89E7F85",
x"A8FA7FB3",
x"A93B7FD0",
x"A96A7FE0",
x"A9917FE8",
x"A9BC7FED",
x"A9F47FF2",
x"AA437FFC",
x"AAB18012",
x"AB438035",
x"ABFA8067",
x"ACD480A9",
x"ADC680F8",
x"AEC98151",
x"AFCA81AC",
x"B0B98202",
x"B185824D",
x"B21E8287",
x"B27E82AB",
x"B2A382BD",
x"B29882C2",
x"B26D82C5",
x"B23D82CF",
x"B22382F1",
x"B2428336",
x"B2AF83A9",
x"B37E844C",
x"B4B6851F",
x"B650861C",
x"B8378735",
x"BA4E8859",
x"BC6E8979",
x"BE6D8A81",
x"C0268B63",
x"C17A8C14",
x"C2578C8A",
x"C2B78CC5",
x"C2A38CC8",
x"C2328C98",
x"C1818C43",
x"C0B28BD3",
x"BFE88B58",
x"BF3F8ADF",
x"BECA8A74",
x"BE918A21",
x"BE8B89E6",
x"BEAA89C5",
x"BED189B4",
x"BEE389A5",
x"BEBF898B",
x"BE4A8955",
x"BD7588F3",
x"BC3C885D",
x"BAA68794",
x"B8CD869C",
x"B6CF8585",
x"B4D48467",
x"B308835C",
x"B1918280",
x"B08B81E8",
x"B00481A5",
x"AFFE81BB",
x"B069821F",
x"B12582C2",
x"B20C8384",
x"B2F18447",
x"B3A884EC",
x"B40B8554",
x"B3FF8571",
x"B377853B",
x"B27184B6",
x"B0F883F0",
x"AF2182FA",
x"AD0481E8",
x"AAB280CC",
x"A83F7FAC",
x"A5B37E88",
x"A30C7D53",
x"A0427BF9",
x"9D457A65",
x"9A03787F",
x"966D7639",
x"92817390",
x"8E42708F",
x"89C36D4E",
x"852769F7",
x"809366BA",
x"7C3963C8",
x"784C6152",
x"74F65F78",
x"72595E56",
x"708C5DEC",
x"6F915E2C",
x"6F605EFD",
x"6FDF6035",
x"70F061A9",
x"726C6334",
x"742F64AF",
x"761D6607",
x"781D672D",
x"7A236824",
x"7C2E68F5",
x"7E4469AE",
x"806C6A62",
x"82B26B1C",
x"851E6BE6",
x"87B16CC5",
x"8A646DB4",
x"8D2C6EAB",
x"8FF76FA4",
x"92AC7094",
x"953B7175",
x"978E7244",
x"999E7302",
x"9B6373B3",
x"9CE3745C",
x"9E277502",
x"9F3E75A7",
x"A032764B",
x"A11276EA",
x"A1E4777E",
x"A2AC77FF",
x"A3667868",
x"A40C78B6",
x"A49B78E7",
x"A50D7901",
x"A566790F",
x"A5AE791D",
x"A5F3793A",
x"A64A796F",
x"A6CA79C9",
x"A7887A46",
x"A8977AE5",
x"A9FD7BA0",
x"ABBB7C68",
x"ADC47D30",
x"B00B7DEB",
x"B2717E91",
x"B4DE7F19",
x"B7387F8B",
x"B9667FE8",
x"BB5B803F",
x"BD0F809B",
x"BE7F810B",
x"BFAF8198",
x"C0A38247",
x"C1648319",
x"C1F58408",
x"C25B8507",
x"C2968605",
x"C2A886F3",
x"C28E87C0",
x"C24A8863",
x"C1E188D0",
x"C1568908",
x"C0B0890D",
x"BFFA88E4",
x"BF39889A",
x"BE788836",
x"BDB987C6",
x"BD018752",
x"BC5086DE",
x"BBA3866D",
x"BAFB85FE",
x"BA538591",
x"B9AC851E",
x"B90284A5",
x"B85B8423",
x"B7BA8399",
x"B726830C",
x"B6A58284",
x"B640820A",
x"B60181A9",
x"B5E9816D",
x"B5FB815D",
x"B633817D",
x"B68881C7",
x"B6E88235",
x"B73C82B1",
x"B76B8328",
x"B75A8382",
x"B6F083A8",
x"B61F838A",
x"B4E1831C",
x"B3428264",
x"B15A816D",
x"AF4F804D",
x"AD507F25",
x"AB917E19",
x"AA3B7D43",
x"A9717CC0",
x"A9457C99",
x"A9AB7CCD",
x"AA8B7D4A",
x"ABB57DF4",
x"ACEE7EA3",
x"ADFD7F30",
x"AEAE7F7A",
x"AEDA7F64",
x"AE747EE5",
x"AD827DFF",
x"AC227CC9",
x"AA7B7B60",
x"A8C079EB",
x"A71C7890",
x"A5B1776B",
x"A487768F",
x"A39875FC",
x"A2C375A3",
x"A1DC7568",
x"A0AE7526",
x"9F0774B1",
x"9CC373EB",
x"99D272B6",
x"9639710C",
x"92186EF5",
x"8DA26C8D",
x"891A69FF",
x"84C6677A",
x"80ED6534",
x"7DC66359",
x"7B7A620E",
x"7A176169",
x"799D6169",
x"79F26201",
x"7AEF6314",
x"7C65647A",
x"7E206609",
x"7FF26797",
x"81B26904",
x"83486A38",
x"84A46B2A",
x"85C86BDC",
x"86BF6C61",
x"87A26CCE",
x"888E6D3F",
x"89A16DCF",
x"8AFA6E96",
x"8CB46FA4",
x"8EDF70FF",
x"918472A6",
x"94A1748D",
x"982876A6",
x"9C0378DA",
x"A0117B12",
x"A4317D3C",
x"A83A7F3F",
x"AC0A8111",
x"AF7882A5",
x"B26E83F3",
x"B4DA84F8",
x"B6AF85B6",
x"B7F0862F",
x"B8A6866A",
x"B8E38670",
x"B8BC864C",
x"B84A860B",
x"B7A885B8",
x"B6EB8560",
x"B628850B",
x"B56E84BF",
x"B4CC847D",
x"B44C8442",
x"B3F7840A",
x"B3D983CC",
x"B3FB8385",
x"B4688331",
x"B52982CF",
x"B6468264",
x"B7BA8200",
x"B98181AC",
x"BB85817E",
x"BDA98184",
x"BFCC81C9",
x"C1C08254",
x"C35E8325",
x"C485842F",
x"C51C8562",
x"C51986A5",
x"C48687DF",
x"C37B88F3",
x"C21B89CC",
x"C08E8A58",
x"BEFF8A87",
x"BD958A5A",
x"BC6489D5",
x"BB788901",
x"BACD87F1",
x"BA5186BC",
x"B9ED8577",
x"B984843B",
x"B8FE831E",
x"B84F8235",
x"B772818B",
x"B674812B",
x"B5678116",
x"B46B8147",
x"B3A381B5",
x"B32C824F",
x"B3218301",
x"B38C83B9",
x"B4708460",
x"B5BC84E4",
x"B7518538",
x"B90A8550",
x"BAB3852B",
x"BC1E84C6",
x"BD188429",
x"BD7D835C",
x"BD35826B",
x"BC388167",
x"BA8C8060",
x"B8517F64",
x"B5AF7E88",
x"B2D97DD6",
x"B0087D57",
x"AD707D14",
x"AB427D0C",
x"A99B7D3A",
x"A8887D95",
x"A8087E0B",
x"A8027E8B",
x"A8537EFE",
x"A8CC7F53",
x"A93D7F78",
x"A97D7F65",
x"A9647F14",
x"A8E17E87",
x"A7F07DC7",
x"A69B7CE5",
x"A4FE7BF4",
x"A3397B04",
x"A1717A25",
x"9FC67962",
x"9E5078C0",
x"9D147837",
x"9C0A77BD",
x"9B1A773D",
x"9A1A769B",
x"98DF75BE",
x"97337490",
x"94F072FB",
x"91F670F6",
x"8E396E85",
x"89C36BB4",
x"84B6689D",
x"7F456563",
x"79B1622F",
x"74425F2E",
x"6F445C87",
x"6AF55A5F",
x"678758CD",
x"651957DF",
x"63B15794",
x"634457DD",
x"63B158A5",
x"64CE59CA",
x"66625B2B",
x"683B5CA1",
x"6A275E0D",
x"6BFD5F56",
x"6DA46069",
x"6F0C6141",
x"703461DD",
x"71246249",
x"71EC6293",
x"72A362CE",
x"735C6309",
x"74286356",
x"751463BF",
x"76256446",
x"775964EC",
x"78A465A8",
x"79FA6670",
x"7B4C673A",
x"7C8967F5",
x"7DA3689B",
x"7E906927",
x"7F4C6994",
x"7FDB69E6",
x"80416A21",
x"80876A4B",
x"80BC6A6B",
x"80EA6A87",
x"811D6AA1",
x"81596ABD",
x"81A56AD5",
x"81FE6AE8",
x"82636AF2",
x"82CC6AED",
x"83376AD9",
x"839A6AB4",
x"83F46A82",
x"84456A47",
x"848B6A0A",
x"84CE69D6",
x"851369B2",
x"856269A7",
x"85C669BA",
x"864669EF",
x"86EC6A45",
x"87B76ABB",
x"88AA6B48",
x"89BE6BE8",
x"8AEC6C8F",
x"8C246D35",
x"8D596DD2",
x"8E776E61",
x"8F706EDC",
x"90326F40",
x"90B66F8C",
x"90F96FBD",
x"90FB6FD5",
x"90C86FD2",
x"906D6FB7",
x"8FFD6F85",
x"8F886F3D",
x"8F226EE5",
x"8ED66E85",
x"8EAB6E26",
x"8EA26DD5",
x"8EBB6D9D",
x"8EEC6D88",
x"8F2B6DA0",
x"8F6E6DE6",
x"8FAE6E5C",
x"8FE46EF9",
x"900E6FAE",
x"902E706F",
x"90427124",
x"904C71BE",
x"904F722B",
x"90487262",
x"9032725A",
x"90077212",
x"8FBE7193",
x"8F5070E6",
x"8EB8701A",
x"8DF16F3D",
x"8CFD6E5E",
x"8BE06D8A",
x"8A9F6CCD",
x"89466C2B",
x"87E06BAA",
x"86776B48",
x"85156B04",
x"83C46AD9",
x"828B6AC2",
x"81746ABA",
x"80896ABE",
x"7FD26AC8",
x"7F5B6AD8",
x"7F2E6AEC",
x"7F556B02",
x"7FD56B1C",
x"80AE6B38",
x"81DC6B55",
x"834F6B73",
x"84F76B92",
x"86B96BAD",
x"887E6BC5",
x"8A2B6BDC",
x"8BA86BF0",
x"8CE26C03",
x"8DCB6C16",
x"8E576C2A",
x"8E866C3A",
x"8E506C42",
x"8DB56C3B",
x"8CAE6C19",
x"8B396BCE",
x"89506B4C",
x"86F06A8C",
x"841B6984",
x"80DD6838",
x"7D4866B0",
x"797C64FA",
x"75A0632F",
x"71E8616D",
x"6E835FD0",
x"6BA75E76",
x"69775D70",
x"68135CCF",
x"67835C95",
x"67BF5CB8",
x"68B15D29",
x"6A325DD3",
x"6C165E9A",
x"6E2D5F67",
x"70486027",
x"724860CE",
x"74106156",
x"759661C3",
x"76D9621F",
x"77E36277",
x"78C562DA",
x"798E6355",
x"7A5563EF",
x"7B2564AA",
x"7C0E6586",
x"7D136677",
x"7E356773",
x"7F73686D",
x"80C76955",
x"82286A21",
x"83906AC8",
x"84F16B47",
x"86456B9D",
x"87836BCF",
x"88A16BE6",
x"899D6BEC",
x"8A716BEB",
x"8B1F6BE9",
x"8BA86BF2",
x"8C136C07",
x"8C656C30",
x"8CA86C68",
x"8CE56CAE",
x"8D246D03",
x"8D6D6D61",
x"8DC56DC5",
x"8E316E33",
x"8EB56EAA",
x"8F566F30",
x"90176FC5",
x"90FD7072",
x"920D7137",
x"93467213",
x"94AA7305",
x"96357400",
x"97DD74FC",
x"999875EC",
x"9B5276C3",
x"9CF87775",
x"9E7A77FF",
x"9FC3785E",
x"A0CC7898",
x"A18B78B6",
x"A20578C7",
x"A24278D8",
x"A24D78F4",
x"A2387922",
x"A2147962",
x"A1ED79B3",
x"A1D07A08",
x"A1BF7A53",
x"A1BB7A86",
x"A1BF7A99",
x"A1C67A84",
x"A1CC7A49",
x"A1CA79F1",
x"A1C07989",
x"A1B37926",
x"A1A878DA",
x"A1A878B4",
x"A1BC78BE",
x"A1EB78FC",
x"A2387964",
x"A29E79EB",
x"A3157A79",
x"A3917AFC",
x"A4007B5E",
x"A44F7B8C",
x"A46E7B7F",
x"A4547B33",
x"A3FB7AAF",
x"A36179FE",
x"A290792F",
x"A18E7850",
x"A06D7771",
x"9F367697",
x"9DF675C8",
x"9CAE7503",
x"9B637441",
x"9A11737F",
x"98B472B6",
x"974971E6",
x"95D07113",
x"94507045",
x"92D26F89",
x"91636EEB",
x"90186E73",
x"8F016E2B",
x"8E286E10",
x"8D916E1D",
x"8D396E43",
x"8D0E6E70",
x"8CFD6E96",
x"8CEC6EA3",
x"8CC26E8F",
x"8C6D6E55",
x"8BE66E00",
x"8B2F6D9C",
x"8A566D3A",
x"89736CEB",
x"889D6CBF",
x"87E76CBB",
x"87606CDC",
x"87066D14",
x"86C56D4B",
x"867E6D65",
x"86096D41",
x"853A6CC4",
x"83E76BD9",
x"81F96A79",
x"7F6368A7",
x"7C356675",
x"78916400",
x"74A8616D",
x"70BA5EE7",
x"6D065C95",
x"69CB5A9B",
x"67355915",
x"65665811",
x"64665794",
x"64305798",
x"64A8580F",
x"65B358E3",
x"672359F8",
x"68D55B38",
x"6AA65C88",
x"6C795DD5",
x"6E3D5F0D",
x"6FE56027",
x"7170611D",
x"72DE61ED",
x"7435629D",
x"757D6332",
x"76C163B7",
x"78076434",
x"795964B2",
x"7ABD653C",
x"7C3565D8",
x"7DC46686",
x"7F606748",
x"81066817",
x"82A568EC",
x"843269BB",
x"859E6A7A",
x"86DD6B1C",
x"87E96B99",
x"88BE6BEC",
x"89626C17",
x"89DD6C1D",
x"8A3E6C0A",
x"8A916BEB",
x"8AE46BCB",
x"8B406BB8",
x"8BA46BBA",
x"8C0A6BD2",
x"8C696C00",
x"8CB16C3E",
x"8CD26C7F",
x"8CC26CB7",
x"8C796CDE",
x"8BFA6CE9",
x"8B4C6CD7",
x"8A806CA8",
x"89A76C66",
x"88D56C1A",
x"881D6BCF",
x"87886B92",
x"871E6B68",
x"86DD6B55",
x"86BE6B59",
x"86B86B6C",
x"86BC6B83",
x"86C56B94",
x"86C86B94",
x"86C36B7C",
x"86B96B48",
x"86AE6AFA",
x"86AA6A9C",
x"86AE6A35",
x"86C369D4",
x"86E76983",
x"871B694E",
x"8759693B",
x"879D694C",
x"87E36980",
x"882769D2",
x"88696A3A",
x"88AB6AB0",
x"88F06B27",
x"893B6B9A",
x"898E6C00",
x"89EA6C55",
x"8A4B6C94",
x"8AA76CBB",
x"8AF46CCA",
x"8B2A6CC1",
x"8B3B6CA3",
x"8B226C75",
x"8ADF6C3E",
x"8A736C06",
x"89E76BD4",
x"894E6BB0",
x"88B26BA0",
x"88276BA6",
x"87B76BBE",
x"87666BE2",
x"87346C09",
x"87186C24",
x"87046C2A",
x"86E66C0C",
x"86AE6BC7",
x"864F6B59",
x"85BF6AC8",
x"85016A20",
x"8421696F",
x"832D68C9",
x"8239683C",
x"815F67D8",
x"80AF67A0",
x"80386794",
x"7FFF67AE",
x"800067E3",
x"80316823",
x"8081685E",
x"80DC6886",
x"812E6894",
x"81686883",
x"81796854",
x"815C680C",
x"810D67B1",
x"808E674C",
x"7FE266E3",
x"7F076676",
x"7E036604",
x"7CD06587",
x"7B7064F7",
x"79DF644E",
x"781B6381",
x"7628628E",
x"74106176",
x"71DC603C",
x"6FA35EEC",
x"6D785D92",
x"6B755C42",
x"69B25B0A",
x"684459FD",
x"67375925",
x"6696588E",
x"6661583F",
x"66965838",
x"672E587A",
x"68235902",
x"696F59D0",
x"6B135AE1",
x"6D105C33",
x"6F6D5DC9",
x"72375FA2",
x"757061BE",
x"79206418",
x"7D4166AE",
x"81C36973",
x"868E6C59",
x"8B7D6F4E",
x"9063723A",
x"95117508",
x"995977A2",
x"9D1479F5",
x"A0227BF5",
x"A2787D98",
x"A4177EDE",
x"A50D7FCA",
x"A574806A",
x"A57180C6",
x"A52880EE",
x"A4BB80EB",
x"A44380C7",
x"A3D28087",
x"A36E8029",
x"A3157FAF",
x"A2B97F14",
x"A24C7E59",
x"A1C07D7A",
x"A10A7C7C",
x"A0247B68",
x"9F117A46",
x"9DDC7923",
x"9C94780F",
x"9B497715",
x"9A10763E",
x"98F77590",
x"9807750C",
x"974674B0",
x"96B27474",
x"96437450",
x"95F1743B",
x"95B37431",
x"9583742F",
x"95607430",
x"954C7439",
x"954D744D",
x"956C746C",
x"95AF749D",
x"961C74DC",
x"96B27529",
x"9764757B",
x"982775CD",
x"98E37616",
x"99837650",
x"99F07677",
x"9A1C7688",
x"9A037685",
x"99A27671",
x"990D7652",
x"9858762F",
x"979D760B",
x"96F875E8",
x"968475C8",
x"964F75AC",
x"96647592",
x"96C1757B",
x"9756756C",
x"9817756A",
x"98ED757E",
x"99C875B3",
x"9A977612",
x"9B5576A0",
x"9BFD7760",
x"9C927848",
x"9D1C794B",
x"9DA17A53",
x"9E247B43",
x"9E9F7BFC",
x"9F117C65",
x"9F697C6A",
x"9F997C01",
x"9F917B2A",
x"9F4379F5",
x"9EA7787C",
x"9DB976DD",
x"9C827539",
x"9B0D73AD",
x"996F7254",
x"97BE7139",
x"96117061",
x"947D6FC3",
x"93156F52",
x"91E06EFA",
x"90E26EA9",
x"90146E4D",
x"8F6C6DD9",
x"8ED66D4B",
x"8E416CA4",
x"8D946BEC",
x"8CBE6B2B",
x"8BAE6A6D",
x"8A5C69BC",
x"88C3691D",
x"86EC6894",
x"84E36820",
x"82BC67BC",
x"808D6768",
x"7E6A671A",
x"7C6966CE",
x"7A93667C",
x"78E9661E",
x"776265AB",
x"75E9651D",
x"74636468",
x"72B16381",
x"70B46262",
x"6E556103",
x"6B8A5F63",
x"685B5D88",
x"64DE5B81",
x"613B5963",
x"5DA75746",
x"5A5B554D",
x"57905396",
x"5575523F",
x"542C515D",
x"53C150FE",
x"54305123",
x"555C51C4",
x"571D52CE",
x"59405426",
x"5B8F55AE",
x"5DDB5745",
x"5FFC58CF",
x"61DC5A35",
x"63725B69",
x"64C15C60",
x"65D85D1B",
x"66CC5DA2",
x"67B55E00",
x"68A75E42",
x"69AE5E76",
x"6ACF5EA8",
x"6C075EE6",
x"6D4F5F35",
x"6E995F98",
x"6FD4600D",
x"70F06093",
x"71E5611D",
x"72A661A5",
x"732E6221",
x"73826287",
x"73A162CF",
x"739662F3",
x"736A62F3",
x"732A62D0",
x"72E26294",
x"729E6246",
x"726B61F2",
x"725261A5",
x"72596168",
x"72866145",
x"72D5613E",
x"73426153",
x"73C96180",
x"745F61BC",
x"74FA61FE",
x"7594623C",
x"76236270",
x"76A56291",
x"7719629F",
x"777D629D",
x"77D6628D",
x"78276276",
x"786D6260",
x"78AD6252",
x"78E0624E",
x"79096258",
x"7920626D",
x"7925628E",
x"791D62B7",
x"790962E2",
x"78F26310",
x"78E6633E",
x"78F0636D",
x"7920639F",
x"797A63D5",
x"7A066413",
x"7ABF6456",
x"7B9E64A3",
x"7C9164F4",
x"7D866546",
x"7E636597",
x"7F1665DF",
x"7F87661B",
x"7FAF6649",
x"7F896666",
x"7F166672",
x"7E636670",
x"7D836665",
x"7C8D6653",
x"7B97663F",
x"7AB7662D",
x"79FF661B",
x"797D660E",
x"79356600",
x"792765F0",
x"794965D9",
x"799065B8",
x"79EA6587",
x"7A476548",
x"7A9464F9",
x"7AC5649B",
x"7ACF6435",
x"7AAB63CE",
x"7A5C6369",
x"79E66310",
x"795162C8",
x"78A76295",
x"77F7627C",
x"774C6279",
x"76B2628D",
x"763162B4",
x"75CE62E4",
x"758C631D",
x"756C6352",
x"7569637F",
x"757F639E",
x"75A763AD",
x"75D963A8",
x"76136390",
x"764C6369",
x"76846337",
x"76BB6301",
x"76F362D2",
x"773062B1",
x"777662A7",
x"77CB62BB",
x"782B62ED",
x"7891633C",
x"78F2639E",
x"79386404",
x"79496459",
x"79066483",
x"784F646A",
x"770963F9",
x"7520631D",
x"728E61D0",
x"6F60601A",
x"6BB55E0B",
x"67BD5BC3",
x"63B4596B",
x"5FE5572E",
x"5C995539",
x"5A1053B5",
x"587F52BD",
x"58055261",
x"58A7529F",
x"5A575368",
x"5CE654A1",
x"60215626",
x"63C157D3",
x"67825984",
x"6B275B1C",
x"6E7C5C8B",
x"71615DC9",
x"73C55ED7",
x"75AA5FBF",
x"771A608E",
x"782E614E",
x"78FA6209",
x"799862C4",
x"7A186379",
x"7A866425",
x"7AE364C1",
x"7B34653F",
x"7B72659D",
x"7B9B65D8",
x"7BAE65F6",
x"7BB165FD",
x"7BA865FA",
x"7B9E65FA",
x"7B9E6604",
x"7BAF6620",
x"7BDC664E",
x"7C236689",
x"7C8366C6",
x"7CF36700",
x"7D6D6728",
x"7DE5673B",
x"7E4F6735",
x"7EA7671A",
x"7EE766F2",
x"7F1466C9",
x"7F2E66AB",
x"7F3F66A4",
x"7F4E66BC",
x"7F6366F7",
x"7F866752",
x"7FBA67C9",
x"80006852",
x"805868E3",
x"80BE6972",
x"812D69F6",
x"81A06A6B",
x"82106ACC",
x"827A6B1C",
x"82D86B57",
x"83256B82",
x"835D6B9C",
x"837D6BA4",
x"83836B9C",
x"836F6B80",
x"83426B54",
x"83036B17",
x"82B86ACC",
x"826F6A7D",
x"82316A30",
x"820B69EF",
x"820A69C4",
x"823569BA",
x"829069D6",
x"83176A19",
x"83C26A7F",
x"84846AFF",
x"85496B8A",
x"85FE6C12",
x"86906C82",
x"86ED6CCD",
x"870D6CE3",
x"86EC6CBF",
x"868A6C63",
x"85F36BD2",
x"85346B1C",
x"845D6A51",
x"837D6986",
x"82A468CE",
x"81D96835",
x"812267C8",
x"80806787",
x"7FEF676D",
x"7F6A6770",
x"7EEC6781",
x"7E706794",
x"7DF56797",
x"7D796783",
x"7D016753",
x"7C8E670B",
x"7C2566AE",
x"7BC66646",
x"7B7365E0",
x"7B256580",
x"7ADB652F",
x"7A8C64EF",
x"7A3464BE",
x"79D16495",
x"79636470",
x"78EF6449",
x"787D641D",
x"781B63E8",
x"77D663AD",
x"77BC6373",
x"77DB6345",
x"783A632B",
x"78DC632F",
x"79BB6359",
x"7ACE63AB",
x"7BFF6424",
x"7D3464BC",
x"7E4B6566",
x"7F256610",
x"7FA266A7",
x"7FA76717",
x"7F22674E",
x"7E0E673E",
x"7C7966E3",
x"7A7C663F",
x"78416560",
x"7601645A",
x"73FD634E",
x"7272625A",
x"719E61A7",
x"71AE6155",
x"72C16180",
x"74DC623C",
x"77F5638D",
x"7BE8656A",
x"808467C4",
x"85916A77",
x"8AD36D63",
x"90147061",
x"9525734A",
x"99E97602",
x"9E4F7875",
x"A2557A9B",
x"A6007C72",
x"A95F7E04",
x"AC827F5D",
x"AF748092",
x"B24381B0",
x"B4F082C3",
x"B77A83D0",
x"B9DA84DC",
x"BC0B85E2",
x"BE0486DC",
x"BFBD87C6",
x"C137889B",
x"C26F895C",
x"C36E8A0A",
x"C43A8AAA",
x"C4DB8B45",
x"C55E8BE0",
x"C5D08C84",
x"C6378D31",
x"C6A28DE9",
x"C7168EA2",
x"C79D8F59",
x"C83F9004",
x"C8FF9098",
x"C9E59116",
x"CAF89179",
x"CC3A91C8",
x"CDB0920E",
x"CF5D9258",
x"D13C92B1",
x"D349932A",
x"D57893C7",
x"D7BD948D",
x"DA069576",
x"DC3D9679",
x"DE519786",
x"E030988F",
x"E1CE9982",
x"E3259A52",
x"E4349AFB",
x"E5039B79",
x"E59C9BCF",
x"E6089C07",
x"E6509C29",
x"E67B9C3D",
x"E6889C47",
x"E6719C4B",
x"E6299C42",
x"E5A79C29",
x"E4E29BF3",
x"E3D89B9C",
x"E2909B1C",
x"E11A9A76",
x"DF9099B0",
x"DE1298D8",
x"DCBE97FD",
x"DBB19735",
x"DAFE9690",
x"DAAD961D",
x"DAB995E3",
x"DB0F95E3",
x"DB989616",
x"DC349670",
x"DCCA96DF",
x"DD3E974F",
x"DD8297B3",
x"DD9097FA",
x"DD68981F",
x"DD12981B",
x"DC9997F2",
x"DC0997AA",
x"DB6A9748",
x"DAC196D9",
x"DA169665",
x"D96795F3",
x"D8B3958D",
x"D7FF9537",
x"D74B94F6",
x"D69D94CF",
x"D5FB94C1",
x"D56B94CF",
x"D4F294F5",
x"D4959531",
x"D453957C",
x"D42995CF",
x"D4169623",
x"D416966E",
x"D42796A7",
x"D44696C8",
x"D46F96CB",
x"D4A596AE",
x"D4E4966E",
x"D5299609",
x"D56F9584",
x"D5B094E3",
x"D5E5942A",
x"D6089360",
x"D6179293",
x"D61391D1",
x"D6029125",
x"D5EB90A2",
x"D5D89053",
x"D5CD903E",
x"D5C19060",
x"D5A390AD",
x"D551910C",
x"D49A9156",
x"D3449165",
x"D1129107",
x"CDC99011",
x"C93E8E60",
x"C3638BE3",
x"BC43889B",
x"B412849F",
x"AB25801C",
x"A1E67B51",
x"98D97688",
x"9080720C",
x"89556E24",
x"83BB6B0A",
x"7FF368E9",
x"7E1A67CF",
x"7E2267BB",
x"7FDD6897",
x"83046A3E",
x"873E6C82",
x"8C2E6F34",
x"91807224",
x"96ED752C",
x"9C407826",
x"A15A7AFE",
x"A62B7D9F",
x"AAAE8000",
x"AEE48219",
x"B2D783ED",
x"B685857A",
x"B9ED86C5",
x"BD0587D6",
x"BFC688B8",
x"C226897A",
x"C4208A2B",
x"C5B68ADA",
x"C6F18B97",
x"C7E18C67",
x"C89D8D50",
x"C93D8E52",
x"C9DD8F63",
x"CA8C9077",
x"CB5E9184",
x"CC54927C",
x"CD6F9356",
x"CEA39410",
x"CFE194AA",
x"D115952B",
x"D22A959B",
x"D30E9603",
x"D3AA9668",
x"D3F696CB",
x"D3E59724",
x"D3749769",
x"D2A2978C",
x"D175977D",
x"CFFF9734",
x"CE5196AD",
x"CC8995EA",
x"CACA9500",
x"C9379403",
x"C7FA9313",
x"C735924C",
x"C70191CB",
x"C77091A0",
x"C88191D1",
x"CA239256",
x"CC36931D",
x"CE889407",
x"D0E294F2",
x"D30995BD",
x"D4CB964E",
x"D5FF9696",
x"D68D9693",
x"D6789652",
x"D5CE95E6",
x"D4B79570",
x"D361950A",
x"D1FF94CE",
x"D0C694CC",
x"CFD8950A",
x"CF53957D",
x"CF3C9614",
x"CF8D96B5",
x"D0339744",
x"D11297A7",
x"D20F97CF",
x"D30F97B5",
x"D3FE9760",
x"D4D396E2",
x"D5899652",
x"D62595CE",
x"D6AA9572",
x"D7259554",
x"D7959582",
x"D7FE95FF",
x"D85B96BF",
x"D8AC97B4",
x"D8E998C4",
x"D91299D1",
x"D9279AC1",
x"D9309B7D",
x"D9399BFB",
x"D9509C30",
x"D9829C21",
x"D9DA9BDC",
x"DA5F9B71",
x"DB0E9AF3",
x"DBDA9A7B",
x"DCB09A17",
x"DD7699D5",
x"DE1099B7",
x"DE6299B8",
x"DE5499CC",
x"DDD599DE",
x"DCDE99D5",
x"DB6C9997",
x"D9899910",
x"D740982D",
x"D4A396E5",
x"D1C3953D",
x"CEB0933F",
x"CB7C9103",
x"C8368EA4",
x"C4EB8C43",
x"C1AB89FE",
x"BE7F87F3",
x"BB758631",
x"B89884BF",
x"B5E98398",
x"B36082A8",
x"B0F081D3",
x"AE7880F2",
x"ABD37FDE",
x"A8C97E70",
x"A5277C82",
x"A0BE7A02",
x"9B6D76EA",
x"95297344",
x"8E076F2B",
x"86366ACE",
x"7E0A6660",
x"75E6621F",
x"6E3F5E48",
x"678C5B10",
x"6230589E",
x"5E78570C",
x"5C89565D",
x"5C625681",
x"5DDB575A",
x"60AA58BD",
x"646B5A78",
x"68B15C59",
x"6D145E36",
x"713B5FEC",
x"74E06166",
x"77DD629D",
x"7A286394",
x"7BCF645A",
x"7CF36500",
x"7DBF659B",
x"7E66663E",
x"7F1066F5",
x"7FDD67C6",
x"80E568B5",
x"822D69BB",
x"83AE6AD1",
x"855C6BE9",
x"871E6CFA",
x"88E06DF8",
x"8A8A6EDC",
x"8C0D6FA3",
x"8D5B7048",
x"8E7070CF",
x"8F53713D",
x"900D7195",
x"90AB71DC",
x"913E721C",
x"91D57254",
x"9279728A",
x"933272BD",
x"940172EC",
x"94DD7317",
x"95BE733B",
x"96927355",
x"97537368",
x"97F47374",
x"9870737C",
x"98CA7386",
x"990B739C",
x"993E73C0",
x"997073F8",
x"99B27447",
x"9A1074AC",
x"9A8D7525",
x"9B2B75AA",
x"9BE67636",
x"9CB576BE",
x"9D8E773E",
x"9E6677AF",
x"9F36780D",
x"9FFA785B",
x"A0B2789B",
x"A16478D1",
x"A21A7908",
x"A2DF794A",
x"A3C279A5",
x"A4CF7A22",
x"A6177AD0",
x"A7A47BBA",
x"A9817CEA",
x"ABB37E64",
x"AE3F8026",
x"B122822C",
x"B4508467",
x"B7B986C2",
x"BB43891F",
x"BECF8B62",
x"C2358D66",
x"C5508F13",
x"C7F89052",
x"CA0E9116",
x"CB7B915D",
x"CC369134",
x"CC4190B1",
x"CBAD8FED",
x"CA998F0B",
x"C9288E28",
x"C7828D60",
x"C5CB8CC3",
x"C4288C5D",
x"C2AC8C2A",
x"C1648C21",
x"C0508C35",
x"BF6A8C50",
x"BE9F8C62",
x"BDE08C58",
x"BD158C27",
x"BC328BC6",
x"BB2F8B38",
x"BA098A7D",
x"B8CD89A1",
x"B78B88B1",
x"B65D87BE",
x"B55D86D9",
x"B4A88617",
x"B4568585",
x"B4778533",
x"B50E8528",
x"B6148563",
x"B77185DC",
x"B9048684",
x"BA9F8745",
x"BC168804",
x"BD3988A5",
x"BDE0890E",
x"BDED8928",
x"BD4E88E7",
x"BC028845",
x"BA0F8742",
x"B78785E7",
x"B47F8443",
x"B10E8260",
x"AD46804D",
x"A93B7E14",
x"A4F07BBA",
x"A0747948",
x"9BCF76C3",
x"970E7436",
x"924C71AF",
x"8DA56F43",
x"89466D0C",
x"855B6B26",
x"821569AA",
x"7FA068AE",
x"7E1B683C",
x"7D956855",
x"7E0B68EB",
x"7F6369E6",
x"81726B26",
x"84006C89",
x"86D36DEF",
x"89B26F41",
x"8C6C7073",
x"8EE07186",
x"91047285",
x"92DF7380",
x"94847490",
x"961875C7",
x"97C27733",
x"99A778D7",
x"9BE67AAC",
x"9E8E7CA2",
x"A1A57EA5",
x"A51E8099",
x"A8DD826B",
x"ACC08407",
x"B09C8563",
x"B447867A",
x"B79C874F",
x"BA7887ED",
x"BCC7885F",
x"BE7F88B2",
x"BFA588F3",
x"C043892B",
x"C0748963",
x"C05489A1",
x"C00989E9",
x"BFB58A3C",
x"BF778A9E",
x"BF6B8B0D",
x"BFA58B8A",
x"C02B8C11",
x"C0FB8C9D",
x"C20B8D27",
x"C3438DA8",
x"C48B8E18",
x"C5C78E71",
x"C6E08EB1",
x"C7C18ED6",
x"C8628EE6",
x"C8C48EE5",
x"C8F48EDD",
x"C9098EDB",
x"C9208EE2",
x"C95B8EFA",
x"C9D88F28",
x"CAB08F69",
x"CBEE8FB9",
x"CD959014",
x"CF939073",
x"D1D190D1",
x"D429912D",
x"D6749187",
x"D88991E2",
x"DA4A9242",
x"DBA092AA",
x"DC82931B",
x"DCF49396",
x"DD059410",
x"DCCD9482",
x"DC6194D8",
x"DBD89504",
x"DB3E94F3",
x"DA989497",
x"D9DE93E6",
x"D90392DE",
x"D7F49184",
x"D69F8FEA",
x"D4FB8E24",
x"D3088C4F",
x"D0D08A87",
x"CE6E88E9",
x"CC02878A",
x"C9B08678",
x"C79D85BF",
x"C5E38556",
x"C48C8535",
x"C3968548",
x"C2ED857A",
x"C26A85B5",
x"C1E385E0",
x"C12685EC",
x"C00B85C8",
x"BE70856C",
x"BC4784D4",
x"B9928402",
x"B66582FB",
x"B2E681C6",
x"AF408070",
x"ABAB7F05",
x"A8547D96",
x"A56A7C32",
x"A30A7AE8",
x"A14879C9",
x"A02278E4",
x"9F8E783E",
x"9F7177E1",
x"9FA877C4",
x"A00A77DE",
x"A069781C",
x"A09F7867",
x"A08B78A2",
x"A01278B6",
x"9F29788B",
x"9DCF7812",
x"9C0E7747",
x"99FE7630",
x"97BE74DB",
x"956C735F",
x"932871DA",
x"910B7061",
x"8F256F0C",
x"8D796DE6",
x"8BFB6CF3",
x"8A976C2A",
x"892E6B78",
x"879E6AC7",
x"85CB69FD",
x"839F690A",
x"811467E0",
x"7E35667F",
x"7B1E64F3",
x"77F76355",
x"74F761BF",
x"72536058",
x"70415F39",
x"6EE65E7E",
x"6E5C5E35",
x"6EA45E5C",
x"6FB05EE9",
x"715F5FC8",
x"738460DD",
x"75F0620D",
x"7873633E",
x"7AE2645D",
x"7D216560",
x"7F246649",
x"80E9671B",
x"827C67E5",
x"83EC68B2",
x"85506993",
x"86BC6A8D",
x"883C6BA4",
x"89D86CD4",
x"8B876E12",
x"8D426F4F",
x"8EF4707E",
x"908D718D",
x"91F77274",
x"9324732A",
x"940E73B3",
x"94B47412",
x"951F7451",
x"95637480",
x"959874B0",
x"95D974EC",
x"96427541",
x"96EC75B7",
x"97E77651",
x"993E770B",
x"9AF077DD",
x"9CF378BD",
x"9F33799C",
x"A1987A71",
x"A4027B30",
x"A6577BD6",
x"A87B7C5E",
x"AA5C7CCE",
x"ABEB7D2D",
x"AD287D87",
x"AE177DE3",
x"AEBF7E49",
x"AF307EBF",
x"AF787F43",
x"AFA57FD6",
x"AFC08070",
x"AFD08108",
x"AFDB8195",
x"AFE48212",
x"AFEA8278",
x"AFF382C6",
x"B00082FD",
x"B01B8322",
x"B04C8339",
x"B09B8347",
x"B1128354",
x"B1B68364",
x"B287837A",
x"B37F8398",
x"B49883C3",
x"B5BF83FE",
x"B6E5844F",
x"B7F884B8",
x"B8E7853D",
x"B9A585DE",
x"BA2B869B",
x"BA75876D",
x"BA8C8849",
x"BA748927",
x"BA3989F4",
x"B9E88AA8",
x"B98C8B35",
x"B92F8B98",
x"B8D48BCD",
x"B8828BDC",
x"B8378BCD",
x"B7F48BAC",
x"B7B98B85",
x"B7858B63",
x"B75E8B4C",
x"B7468B3F",
x"B7468B39",
x"B7618B31",
x"B79B8B17",
x"B7F48ADF",
x"B8638A7D",
x"B8DB89E9",
x"B94C891E",
x"B99C881F",
x"B9B586F8",
x"B98185B5",
x"B8F4846A",
x"B80B832C",
x"B6CF820F",
x"B5568129",
x"B3C08087",
x"B2358030",
x"B0DD802C",
x"AFDD8071",
x"AF4D80F4",
x"AF3C81A3",
x"AFA28267",
x"B06B8326",
x"B17783CC",
x"B29F8447",
x"B3BA848E",
x"B4AB849F",
x"B5578485",
x"B5B98450",
x"B5D48414",
x"B5B683E4",
x"B56E83D2",
x"B50883E1",
x"B485840A",
x"B3D78436",
x"B2E08445",
x"B1708408",
x"AF538357",
x"AC568207",
x"A84F7FFC",
x"A32B7D32",
x"9CF879AF",
x"95E77599",
x"8E457129",
x"867C6CA4",
x"7F036856",
x"78526489",
x"72D86176",
x"6EE05F48",
x"6C9B5E14",
x"6C0D5DD3",
x"6D0D5E6C",
x"6F595FB1",
x"7291616D",
x"764C6368",
x"7A27656A",
x"7DC9674B",
x"80F068E8",
x"83796A30",
x"85586B21",
x"869B6BC1",
x"87656C20",
x"87DC6C4E",
x"882B6C62",
x"88766C6B",
x"88D66C76",
x"895A6C8F",
x"8A006CB7",
x"8ABF6CF0",
x"8B896D3A",
x"8C4B6D8F",
x"8CF96DEC",
x"8D876E4D",
x"8DF46EB0",
x"8E426F10",
x"8E776F70",
x"8E9D6FCD",
x"8EB77026",
x"8EC97078",
x"8ED370C0",
x"8ECC70FB",
x"8EAA7120",
x"8E637129",
x"8DED710F",
x"8D4370CB",
x"8C69705B",
x"8B666FC0",
x"8A496EFE",
x"89286E1E",
x"881B6D31",
x"87396C47",
x"86986B73",
x"86436AC7",
x"86456A4F",
x"869B6A1A",
x"873E6A2B",
x"88216A7F",
x"89346B10",
x"8A646BD4",
x"8BA46CBD",
x"8CDF6DBA",
x"8E0D6EBF",
x"8F226FC0",
x"901A70B1",
x"90EC718A",
x"91957244",
x"921472D5",
x"9264733A",
x"9284736A",
x"9274735E",
x"92327315",
x"91C0728C",
x"912571C7",
x"906370D2",
x"8F846FBD",
x"8E926E99",
x"8D9B6D7F",
x"8CAA6C82",
x"8BCF6BB8",
x"8B176B2D",
x"8A906AE3",
x"8A436ADC",
x"8A376B09",
x"8A6C6B59",
x"8ADD6BBA",
x"8B836C19",
x"8C4C6C68",
x"8D246C9E",
x"8DF76CBD",
x"8EB16CCA",
x"8F416CD1",
x"8F986CE2",
x"8FB26D09",
x"8F946D4F",
x"8F426DB7",
x"8ECB6E3B",
x"8E3E6ECF",
x"8DAE6F64",
x"8D256FE4",
x"8CAE7040",
x"8C4F706C",
x"8C097066",
x"8BD57031",
x"8BAE6FD9",
x"8B906F70",
x"8B746F0D",
x"8B5A6EC1",
x"8B426E9D",
x"8B2E6EAA",
x"8B216EE8",
x"8B216F51",
x"8B316FD8",
x"8B4F7069",
x"8B7B70F2",
x"8BB17164",
x"8BE971AF",
x"8C1D71CD",
x"8C4671BD",
x"8C607180",
x"8C63711D",
x"8C48709D",
x"8C077002",
x"8B956F52",
x"8AE46E8C",
x"89E66DAB",
x"88866CAB",
x"86B96B86",
x"84746A35",
x"81B868BC",
x"7E90671E",
x"7B136565",
x"7762639F",
x"73AE61E0",
x"7026603E",
x"6CFD5EC8",
x"6A615D90",
x"68735CA2",
x"674A5C06",
x"66E85BBD",
x"67425BC3",
x"68445C12",
x"69CA5CA1",
x"6BAD5D63",
x"6DCB5E4F",
x"6FFF5F5A",
x"7230607A",
x"744B61A7",
x"764462D9",
x"781B6409",
x"79D2652F",
x"7B726649",
x"7D006753",
x"7E89684B",
x"80116931",
x"81A16A06",
x"833B6ACE",
x"84DF6B8A",
x"86886C3E",
x"88376CE8",
x"89E06D89",
x"8B7F6E1D",
x"8D0A6EA1",
x"8E796F13",
x"8FC56F70",
x"90E76FB9",
x"91DA6FEC",
x"929B7013",
x"93287033",
x"93817051",
x"93A87078",
x"93A170AD",
x"937070F4",
x"931D714D",
x"92B171B9",
x"92397231",
x"91C272B7",
x"915D7344",
x"911B73D7",
x"910B746E",
x"913B7508",
x"91B475A5",
x"92747644",
x"937976E2",
x"94B2777B",
x"960B7806",
x"976C787C",
x"98B978D6",
x"99E07908",
x"9ACD7913",
x"9B7D78F8",
x"9BEE78B9",
x"9C2F7862",
x"9C557801",
x"9C7477A0",
x"9CA57751",
x"9CFA771B",
x"9D7E7705",
x"9E32770D",
x"9F0D7731",
x"9FFE7765",
x"A0F0779F",
x"A1CD77D0",
x"A28177F1",
x"A2FE77F9",
x"A33B77EA",
x"A33C77C3",
x"A308778D",
x"A2B17752",
x"A246771C",
x"A1D976F2",
x"A17776DD",
x"A12876DD",
x"A0ED76F4",
x"A0C37719",
x"A0A17747",
x"A0777772",
x"A03C7792",
x"9FE17799",
x"9F607783",
x"9EB1774A",
x"9DD376EC",
x"9CC9766A",
x"9B9875C7",
x"9A467506",
x"98DC7430",
x"975F734B",
x"95D9725E",
x"94527170",
x"92CC7089",
x"914F6FB0",
x"8FDF6EE9",
x"8E836E3E",
x"8D3F6DB1",
x"8C186D45",
x"8B146CFF",
x"8A356CD9",
x"897D6CD4",
x"88EC6CE6",
x"887D6D09",
x"88286D2E",
x"87E76D4D",
x"87AE6D58",
x"87736D4B",
x"872B6D20",
x"86D16CD7",
x"865C6C73",
x"85CE6C02",
x"85286B8C",
x"84706B1C",
x"83AB6ABA",
x"82DC6A6F",
x"82046A35",
x"81256A0A",
x"803869DF",
x"7F3569A3",
x"7E146944",
x"7CCE68B0",
x"7B5B67D9",
x"79C166BF",
x"78076565",
x"763E63D8",
x"747C622F",
x"72DE608A",
x"717D5F07",
x"70735DCB",
x"6FD55CEE",
x"6FAA5C87",
x"6FF55C9F",
x"70AA5D35",
x"71BA5E3B",
x"730D5F9D",
x"748C613C",
x"762062FC",
x"77B764BB",
x"79456662",
x"7AC967DB",
x"7C45691B",
x"7DC46A26",
x"7F4F6AFF",
x"80F46BB5",
x"82BE6C5B",
x"84B26D00",
x"86D26DB5",
x"89186E83",
x"8B7D6F6B",
x"8DF07066",
x"9063716C",
x"92C3726A",
x"95017350",
x"970B740B",
x"98D87490",
x"9A5C74DA",
x"9B9474EA",
x"9C8174CA",
x"9D247489",
x"9D84743A",
x"9DAE73F1",
x"9DAC73BE",
x"9D8E73AF",
x"9D6273C8",
x"9D35740B",
x"9D18746E",
x"9D1474EA",
x"9D327571",
x"9D7875F8",
x"9DED7678",
x"9E8D76EC",
x"9F597755",
x"A04A77BA",
x"A15C7822",
x"A2857896",
x"A3BD791D",
x"A4FB79BE",
x"A6337A79",
x"A75A7B49",
x"A8677C28",
x"A9507D09",
x"AA117DE4",
x"AA9F7EAA",
x"AAFB7F53",
x"AB227FD9",
x"AB178035",
x"AADC8066",
x"AA77806D",
x"A9F1804A",
x"A9538004",
x"A8A87F9C",
x"A7FD7F19",
x"A75E7E7F",
x"A6D77DD4",
x"A6757D20",
x"A6407C6B",
x"A63F7BBF",
x"A6757B25",
x"A6E17AA6",
x"A77D7A4A",
x"A83D7A19",
x"A9187A13",
x"A9FD7A3C",
x"AADD7A8B",
x"ABA97AFE",
x"AC577B89",
x"ACDE7C26",
x"AD3D7CC9",
x"AD777D68",
x"AD917E01",
x"AD947E8C",
x"AD897F08",
x"AD7A7F78",
x"AD707FDB",
x"AD6B8033",
x"AD6B8080",
x"AD6A80BC",
x"AD5A80E6",
x"AD2C80F0",
x"ACCF80D4",
x"AC308085",
x"AB457FFE",
x"AA057F39",
x"A8747E3A",
x"A69C7D08",
x"A4927BB2",
x"A2737A4B",
x"A05D78EE",
x"9E7177AF",
x"9CCC76A3",
x"9B8175D7",
x"9A977550",
x"9A087508",
x"99C274F2",
x"99A474FB",
x"99877506",
x"99457501",
x"98B974D1",
x"97CA746A",
x"966E73C6",
x"94AA72E8",
x"929071DC",
x"904270B3",
x"8DE76F7E",
x"8BAA6E51",
x"89A76D3A",
x"87F46C3F",
x"86976B63",
x"85806A9D",
x"849069DE",
x"839B6913",
x"8274682A",
x"80ED6713",
x"7EE665C1",
x"7C4F6434",
x"792E6270",
x"759E6086",
x"71D25E8E",
x"6E095CA7",
x"6A875AEB",
x"67945980",
x"65685877",
x"642A57E7",
x"63E957D4",
x"649C5839",
x"66245908",
x"684E5A2B",
x"6ADC5B81",
x"6D905CEC",
x"702E5E4B",
x"72875F87",
x"747F608D",
x"76096153",
x"772B61D8",
x"77FD6224",
x"789B6246",
x"79286252",
x"79C2625C",
x"7A846277",
x"7B7A62B4",
x"7CAA631D",
x"7E0A63B7",
x"7F8E647F",
x"8121656D",
x"82AD6677",
x"841B678E",
x"856068A6",
x"867169AE",
x"874C6AA0",
x"87F46B76",
x"88746C2D",
x"88D86CC8",
x"892F6D4F",
x"898A6DC7",
x"89F36E38",
x"8A746EA6",
x"8B136F14",
x"8BCE6F82",
x"8CA46FEC",
x"8D8E704E",
x"8E8470A4",
x"8F8070E9",
x"907C7120",
x"9173714A",
x"9266716F",
x"9356719A",
x"944B71D8",
x"95497233",
x"965672B6",
x"97787365",
x"98B4743E",
x"9A04753E",
x"9B677658",
x"9CD3777B",
x"9E3C7895",
x"9F957992",
x"A0CF7A65",
x"A1DC7AFF",
x"A2B27B5D",
x"A3497B78",
x"A3A17B57",
x"A3B97AFF",
x"A39A7A7C",
x"A34B79D7",
x"A2D7791F",
x"A24D785D",
x"A1B9779F",
x"A12276EC",
x"A0957651",
x"A01575D5",
x"9FA97581",
x"9F53755A",
x"9F177562",
x"9EF4759F",
x"9EEE7609",
x"9F04769D",
x"9F357750",
x"9F807810",
x"9FDD78D4",
x"A0487986",
x"A0B67A1C",
x"A11F7A8B",
x"A17A7ACB",
x"A1BF7AE1",
x"A1EA7AD1",
x"A1FA7AA9",
x"A1EE7A72",
x"A1CD7A3E",
x"A19C7A16",
x"A1607A01",
x"A11A79FC",
x"A0C87A03",
x"A0647A06",
x"9FE479F5",
x"9F3E79C0",
x"9E647956",
x"9D4F78B2",
x"9BFB77D0",
x"9A6D76BC",
x"98B47585",
x"96E07444",
x"950B7315",
x"93507210",
x"91C3714D",
x"907670DA",
x"8F7270B7",
x"8EB570DF",
x"8E357140",
x"8DE071C3",
x"8DA5724A",
x"8D6D72BD",
x"8D2B7303",
x"8CD37310",
x"8C6372DC",
x"8BE0726B",
x"8B4F71C1",
x"8AB970EF",
x"8A247005",
x"898B6F0F",
x"88EA6E1A",
x"882D6D2A",
x"873C6C41",
x"86006B59",
x"845C6A6D",
x"82426972",
x"7FAA685E",
x"7C9A672D",
x"792865D9",
x"757D6466",
x"71C862DC",
x"6E3E6146",
x"6B175FB2",
x"68865E33",
x"66B05CDA",
x"65AB5BBB",
x"657D5AE0",
x"661C5A57",
x"676C5A28",
x"694B5A52",
x"6B925AD3",
x"6E135BA4",
x"70AD5CB6",
x"73445DFD",
x"75C45F67",
x"782660E4",
x"7A686263",
x"7C9163D6",
x"7EAC6532",
x"80C3666F",
x"82DF678A",
x"85046883",
x"8734695F",
x"896C6A28",
x"8BA46AE9",
x"8DD56BAD",
x"8FF36C80",
x"91F96D6E",
x"93DF6E7C",
x"959E6FAB",
x"973570FC",
x"98A27265",
x"99E773D8",
x"9B04754A",
x"9BF876A5",
x"9CC777DD",
x"9D6E78E5",
x"9DF079B4",
x"9E4C7A4B",
x"9E887AAD",
x"9EA87AE4",
x"9EB67AFC",
x"9EBD7B02",
x"9ECD7B04",
x"9EF37B0B",
x"9F3E7B1C",
x"9FBB7B3A",
x"A0717B64",
x"A1667B98",
x"A2947BD1",
x"A3F07C0E",
x"A56C7C50",
x"A6F47C99",
x"A8737CED",
x"A9D47D51",
x"AB0C7DC9",
x"AC0F7E54",
x"ACDE7EF1",
x"AD7B7F96",
x"ADF7803D",
x"AE5E80D6",
x"AEC08156",
x"AF2E81B2",
x"AFAC81E3",
x"B04081EA",
x"B0E681CA",
x"B192818E",
x"B23D8143",
x"B2D980FB",
x"B35E80C3",
x"B3C980AC",
x"B42180BD",
x"B46D80FD",
x"B4C2816B",
x"B5308202",
x"B5CA82BC",
x"B69F8388",
x"B7B2845D",
x"B901852E",
x"BA7A85ED",
x"BC078692",
x"BD898719",
x"BEE18781",
x"BFF187C8",
x"C09F87F1",
x"C0DD8803",
x"C0A68803",
x"C00287F6",
x"BEFF87E0",
x"BDB687C5",
x"BC4087A5",
x"BAB6877D",
x"B933874A",
x"B7C7870A",
x"B67E86B9",
x"B55E8656",
x"B46685E0",
x"B392855A",
x"B2DC84CA",
x"B23D8439",
x"B1AF83AD",
x"B12D8332",
x"B0B282CC",
x"B039827D",
x"AFB98246",
x"AF29821F",
x"AE7E8200",
x"ADAB81DC",
x"ACA581A3",
x"AB5E814D",
x"A9D780CD",
x"A8128023",
x"A61F7F50",
x"A4127E5B",
x"A2077D50",
x"A0187C3C",
x"9E627B2A",
x"9CF17A26",
x"9BCC7930",
x"9AE77846",
x"9A287761",
x"996D7672",
x"988B756E",
x"975A744A",
x"95BB72FF",
x"939C7193",
x"9100700C",
x"8DFD6E7F",
x"8ABB6CFF",
x"87696BA3",
x"84426A80",
x"817969A6",
x"7F376917",
x"7D9868D2",
x"7CA768CE",
x"7C5E68F9",
x"7CAA6944",
x"7D7569A1",
x"7EA56A09",
x"80226A77",
x"81E26AF6",
x"83DA6B8C",
x"860E6C4A",
x"88846D3D",
x"8B426E6F",
x"8E4D6FE5",
x"91A2719D",
x"9536738F",
x"98F975A9",
x"9CCF77DA",
x"A09F7A0C",
x"A4497C2F",
x"A7B37E30",
x"AAC78002",
x"AD7881A2",
x"AFC2830B",
x"B1A5843F",
x"B32D8545",
x"B46D8625",
x"B57886EC",
x"B66487A4",
x"B745885C",
x"B829891A",
x"B91E89E9",
x"BA238AC8",
x"BB368BB5",
x"BC4D8CA8",
x"BD578D97",
x"BE468E73",
x"BF0A8F2E",
x"BF988FBE",
x"BFF2901B",
x"C01E9048",
x"C02B9049",
x"C030902F",
x"C047900C",
x"C08B8FF2",
x"C10F8FF4",
x"C1E09021",
x"C3019080",
x"C4689110",
x"C60691CB",
x"C7C192A1",
x"C97F9382",
x"CB25945B",
x"CC99951A",
x"CDCD95B1",
x"CEB49614",
x"CF4B963F",
x"CF929631",
x"CF8C95EE",
x"CF3C957D",
x"CEA794E9",
x"CDD1943E",
x"CCBF9387",
x"CB7592D2",
x"CA01922E",
x"C87191A8",
x"C6DB914B",
x"C55D9124",
x"C4159137",
x"C31E918A",
x"C292921A",
x"C28192E0",
x"C2ED93D1",
x"C3CA94DC",
x"C50195EE",
x"C66A96F5",
x"C7D897D9",
x"C91C988D",
x"CA089903",
x"CA779930",
x"CA4E9910",
x"C98898A7",
x"C82997F8",
x"C6449709",
x"C3F995E8",
x"C16D949B",
x"BEC1932F",
x"BC1C91AD",
x"B999901B",
x"B74A8E81",
x"B53A8CE6",
x"B36E8B4C",
x"B1E089BB",
x"B0858836",
x"AF5686C6",
x"AE44856E",
x"AD468435",
x"AC53831B",
x"AB618226",
x"AA6D8154",
x"A97580A6",
x"A8788016",
x"A7747F9F",
x"A6677F3C",
x"A5547EE3",
x"A43C7E8A",
x"A3217E2A",
x"A2037DBC",
x"A0E97D3C",
x"9FDA7CA8",
x"9EE47C04",
x"9E147B54",
x"9D767AA5",
x"9D1A7A02",
x"9D0A7979",
x"9D487916",
x"9DC878E0",
x"9E7478D3",
x"9F2278E5",
x"9F9C78FF",
x"9F9E7901",
x"9EE078C3",
x"9D22781B",
x"9A3176E2",
x"95F47501",
x"9076726A",
x"89E36F2A",
x"82906B62",
x"7AED6746",
x"73826321",
x"6CD65F3E",
x"67695BEA",
x"63A35967",
x"61C157E7",
x"61D95781",
x"63D45832",
x"677259E0",
x"6C585C5C",
x"721E5F6A",
x"785862CB",
x"7EA46641",
x"84B8699A",
x"8A606CB1",
x"8F806F73",
x"941271DA",
x"981E73EA",
x"9BAC75B1",
x"9ECA7740",
x"A18078A5",
x"A3CC79ED",
x"A5A97B1C",
x"A7127C34",
x"A8007D33",
x"A8747E12",
x"A87D7ECD",
x"A82F7F5D",
x"A7A87FC3",
x"A70A7FFC",
x"A677800C",
x"A60B7FFA",
x"A5D67FC9",
x"A5DA7F7F",
x"A60E7F25",
x"A65D7EC1",
x"A6AB7E5A",
x"A6DA7DF4",
x"A6D07D91",
x"A67E7D35",
x"A5DC7CE0",
x"A4F37C8F",
x"A3D57C40",
x"A29F7BED",
x"A1737B93",
x"A06E7B2F",
x"9FAE7ABD",
x"9F457A44",
x"9F3B79C6",
x"9F8D794B",
x"A02C78E1",
x"A1077893",
x"A200786B",
x"A2FD7877",
x"A3EA78B6",
x"A4B2792D",
x"A54C79D6",
x"A5B37AA3",
x"A5EE7B86",
x"A6047C6B",
x"A6007D3C",
x"A5EA7DE4",
x"A5CA7E53",
x"A59E7E7A",
x"A5607E51",
x"A5057DD7",
x"A47D7D12",
x"A3BC7C0F",
x"A2B67ADE",
x"A16D7999",
x"9FEA7857",
x"9E407731",
x"9C927641",
x"9B047599",
x"99C07547",
x"98ED7552",
x"98A875BA",
x"99047678",
x"9A01777E",
x"9B9478BD",
x"9DA27A22",
x"A00B7B99",
x"A2A47D11",
x"A5467E7A",
x"A7D27FC7",
x"AA2E80F2",
x"AC4681F2",
x"AE1582C2",
x"AF9C835C",
x"B0DD83BC",
x"B1DD83E0",
x"B2A383C7",
x"B3358376",
x"B39282F1",
x"B3C38246",
x"B3C98187",
x"B3AC80C7",
x"B375801E",
x"B3337FA2",
x"B2F47F67",
x"B2C97F78",
x"B2BF7FDB",
x"B2E4808E",
x"B3428182",
x"B3DC82A6",
x"B4AD83E1",
x"B5B3851C",
x"B6E1863F",
x"B826873B",
x"B9748803",
x"BABA8898",
x"BBED8901",
x"BCFE8949",
x"BDEE8984",
x"BEBC89C5",
x"BF728A1F",
x"C01F8AA4",
x"C0D38B5A",
x"C1998C42",
x"C27A8D55",
x"C36D8E7D",
x"C45B8F9E",
x"C51E9091",
x"C577912D",
x"C5229142",
x"C3D690AA",
x"C1508F43",
x"BD608CFD",
x"B7F189D2",
x"B11685D6",
x"A9078130",
x"A01E7C18",
x"96D576CE",
x"8DB671A0",
x"854C6CD8",
x"7E1068B7",
x"78606570",
x"74746321",
x"725561D3",
x"71E16177",
x"72D561ED",
x"74D56307",
x"777A648D",
x"7A5D6649",
x"7D2B680A",
x"7FA169A6",
x"81A06B03",
x"831A6C14",
x"84226CDB",
x"84D66D61",
x"855F6DB8",
x"85E26DF6",
x"86816E2B",
x"87566E69",
x"88666EB7",
x"89AD6F16",
x"8B186F82",
x"8C916FF0",
x"8DFD7054",
x"8F4170A3",
x"904870D1",
x"910470DA",
x"917170BB",
x"9195707C",
x"917B7023",
x"91356FBA",
x"90D56F4E",
x"906C6EEB",
x"90086E9A",
x"8FB36E5F",
x"8F706E3E",
x"8F376E34",
x"8F006E41",
x"8EBF6E5C",
x"8E666E82",
x"8DEA6EAB",
x"8D486ED7",
x"8C806F00",
x"8B9A6F24",
x"8AA46F43",
x"89B26F5B",
x"88D96F6C",
x"882B6F78",
x"87B86F7C",
x"87876F7A",
x"879D6F75",
x"87F26F68",
x"887A6F59",
x"89286F48",
x"89E96F37",
x"8AAF6F27",
x"8B706F19",
x"8C246F0F",
x"8CCB6F0A",
x"8D656F0D",
x"8DFA6F1A",
x"8E8D6F30",
x"8F226F52",
x"8FB96F82",
x"904F6FBD",
x"90D87003",
x"914B704F",
x"919B709F",
x"91BE70E9",
x"91A87126",
x"9158714E",
x"90CE7158",
x"900E7141",
x"8F247102",
x"8E18709F",
x"8CFA701A",
x"8BD56F7A",
x"8AB56ECA",
x"89A76E13",
x"88B16D62",
x"87DF6CBF",
x"87356C34",
x"86BC6BC5",
x"867A6B76",
x"86706B45",
x"86A26B31",
x"870B6B32",
x"87A86B48",
x"886F6B6C",
x"89526B9C",
x"8A486BD7",
x"8B3F6C1D",
x"8C2C6C72",
x"8D046CD8",
x"8DBF6D51",
x"8E5C6DDE",
x"8EDA6E7C",
x"8F416F26",
x"8F946FD5",
x"8FDD7082",
x"9022711F",
x"906671A6",
x"90AC720F",
x"90F07255",
x"912C7278",
x"91597279",
x"916F725C",
x"91667229",
x"913871E6",
x"90E7719A",
x"9073714A",
x"8FE470F6",
x"8F4170A4",
x"8E907052",
x"8DD76FFC",
x"8D186F9D",
x"8C496F31",
x"8B5C6EB0",
x"8A416E13",
x"88E26D51",
x"872B6C65",
x"85116B4B",
x"82946A07",
x"7FC1689E",
x"7CB56724",
x"79A165AF",
x"76BE6460",
x"744E6358",
x"728D62B7",
x"71B2629B",
x"71E26315",
x"7328642D",
x"757C65D3",
x"78B867F0",
x"7CA76A5C",
x"81036CEB",
x"85866F69",
x"89EA71B0",
x"8DF973A0",
x"918B752C",
x"948E7654",
x"97077729",
x"990B77C6",
x"9ABB784D",
x"9C3F78E1",
x"9DC5799F",
x"9F6E7A9C",
x"A1597BE0",
x"A3957D6A",
x"A6287F2D",
x"A908811F",
x"AC298328",
x"AF718536",
x"B2CC873E",
x"B61C8931",
x"B94C8B0B",
x"BC478CC8",
x"BEFC8E65",
x"C1648FDF",
x"C3729134",
x"C528925F",
x"C681935B",
x"C77E9423",
x"C82094B3",
x"C86D9506",
x"C864951B",
x"C80F94F3",
x"C7729493",
x"C69C93FF",
x"C596933E",
x"C4749258",
x"C3449156",
x"C21B9044",
x"C1028F28",
x"C0058E0A",
x"BF298CF3",
x"BE688BE6",
x"BDBA8AE7",
x"BD1489F4",
x"BC65890F",
x"BBA58835",
x"BACE8766",
x"B9E386A1",
x"B8ED85E7",
x"B801853F",
x"B73084AC",
x"B6918436",
x"B63083E0",
x"B61583AC",
x"B6388398",
x"B687839F",
x"B6E883B8",
x"B73C83D3",
x"B76583E7",
x"B75083E8",
x"B6F383D3",
x"B65683AB",
x"B5948377",
x"B4D1834C",
x"B43C833B",
x"B404835A",
x"B44983BB",
x"B5238464",
x"B68F8556",
x"B8748681",
x"BAA687CC",
x"BCE88915",
x"BEF78A35",
x"C0938B07",
x"C18B8B6F",
x"C1C38B5C",
x"C1378ACC",
x"C00489CF",
x"BE568883",
x"BC6E870F",
x"BA9785A1",
x"B9118463",
x"B8128377",
x"B7B782F4",
x"B80482DD",
x"B8E38326",
x"BA2383B6",
x"BB8B846C",
x"BCDB8521",
x"BDD985B3",
x"BE5A860A",
x"BE4A8619",
x"BDAF85E3",
x"BCA28571",
x"BB4E84DD",
x"B9EB843C",
x"B8A983A8",
x"B7B2832D",
x"B71B82D6",
x"B6E4829C",
x"B6FA8274",
x"B733824A",
x"B763820B",
x"B75981A6",
x"B6EA8114",
x"B5FF8050",
x"B4957F64",
x"B2B97E64",
x"B08C7D5E",
x"AE367C6B",
x"ABE67B99",
x"A9BB7AF4",
x"A7C97A79",
x"A6157A20",
x"A48879D4",
x"A300797F",
x"A14C7901",
x"9F3C7841",
x"9CA77729",
x"997475AC",
x"95A273C6",
x"9149717F",
x"8C956EEE",
x"87CB6C2E",
x"83346969",
x"7F1D66C6",
x"7BC96470",
x"796F628D",
x"782A613B",
x"7800608E",
x"78DF6090",
x"7AA3613C",
x"7D176284",
x"8007644F",
x"8338667C",
x"867D68E9",
x"89AF6B72",
x"8CB66DF5",
x"8F867058",
x"921B7285",
x"947D7471",
x"96B57615",
x"98CF7772",
x"9AD77893",
x"9CD77982",
x"9ED37A4D",
x"A0D07B05",
x"A2D07BB7",
x"A4CF7C71",
x"A6CA7D39",
x"A8BF7E12",
x"AAA67EFC",
x"AC7D7FF0",
x"AE3980E6",
x"AFD781D1",
x"B14F82A9",
x"B2988364",
x"B3AF83FE",
x"B48C847B",
x"B52E84E1",
x"B58F8539",
x"B5B5858F",
x"B59F85EC",
x"B5538654",
x"B4D786C9",
x"B4358742",
x"B37587B3",
x"B2A6880D",
x"B1D0883C",
x"B1008833",
x"B03F87E9",
x"AF92875E",
x"AEFE8699",
x"AE8285AB",
x"AE1784A9",
x"ADB683AC",
x"AD5682C9",
x"ACED8216",
x"AC71819C",
x"ABDD8160",
x"AB35815E",
x"AA7E818B",
x"A9C581DA",
x"A91A823D",
x"A88F82A5",
x"A83A8307",
x"A82C835D",
x"A87183A8",
x"A91283E4",
x"AA0A8417",
x"AB4F8442",
x"ACD28467",
x"AE7A8485",
x"B030849C",
x"B1DC84AC",
x"B36784B5",
x"B4C284B9",
x"B5E484BF",
x"B6D084D0",
x"B78C84F8",
x"B8288546",
x"B8B685C2",
x"B94D8674",
x"B9FF8760",
x"BADD8880",
x"BBF189C9",
x"BD428B2C",
x"BECD8C94",
x"C08E8DF0",
x"C2788F2F",
x"C47E9045",
x"C68E912B",
x"C89391E2",
x"CA7B926F",
x"CC2F92D8",
x"CD989324",
x"CEA29359",
x"CF3A9378",
x"CF53937C",
x"CEE79362",
x"CDFB9324",
x"CCA092BD",
x"CAF1922B",
x"C9139173",
x"C72F909D",
x"C5718FB5",
x"C3FC8ECB",
x"C2EE8DEA",
x"C24D8D1E",
x"C2158C69",
x"C22F8BC9",
x"C2758B38",
x"C2C28AAC",
x"C2E88A1F",
x"C2CA898A",
x"C25388F0",
x"C1818857",
x"C05E87CC",
x"BF05875D",
x"BD918712",
x"BC1C86F1",
x"BAB386F1",
x"B95686FA",
x"B7ED86ED",
x"B65186A2",
x"B44D85EC",
x"B1A984A3",
x"AE3882B1",
x"A9D9800B",
x"A4887CC0",
x"9E6678F4",
x"97AC74DC",
x"90B670BB",
x"89ED6CD8",
x"83C26972",
x"7E9B66BF",
x"7ACC64E0",
x"788963DF",
x"77DD63B2",
x"78B5643C",
x"7AD96552",
x"7DFC66C4",
x"81BF6865",
x"85CB6A0C",
x"89CF6BA1",
x"8D926D17",
x"90F66E6C",
x"93F06FAE",
x"969270EE",
x"98F97240",
x"9B4873B3",
x"9D9F7554",
x"A0127725",
x"A2A4791B",
x"A5467B25",
x"A7DD7D2C",
x"AA437F14",
x"AC5080C3",
x"ADE48222",
x"AEF18323",
x"AF7883BF",
x"AF8F83FB",
x"AF6083E3",
x"AF1B838E",
x"AEFD8317",
x"AF36829B",
x"AFED8235",
x"B13581FE",
x"B30A8208",
x"B551825A",
x"B7E082F7",
x"BA7F83D4",
x"BCF384E4",
x"BF068611",
x"C08F8740",
x"C175885C",
x"C1B3894C",
x"C15889FB",
x"C0828A5C",
x"BF5A8A66",
x"BE128A1A",
x"BCD78980",
x"BBD388A2",
x"BB268798",
x"BAE48678",
x"BB13855E",
x"BBAC8463",
x"BC9E839C",
x"BDCA831E",
x"BF0F82F0",
x"C0478311",
x"C14A8378",
x"C1F48412",
x"C22684C5",
x"C1CC8576",
x"C0DA8605",
x"BF568660",
x"BD518673",
x"BAEA863C",
x"B84D85C0",
x"B5A98511",
x"B3358446",
x"B11E837D",
x"AF8C82D0",
x"AE9B8257",
x"AE538223",
x"AEAE8237",
x"AF96828F",
x"B0EA831C",
x"B27E83CA",
x"B4288481",
x"B5BF8529",
x"B72085AF",
x"B8358607",
x"B8ED8628",
x"B9468612",
x"B94085CA",
x"B8E38559",
x"B83384C5",
x"B7398415",
x"B5F7834F",
x"B4708276",
x"B2A6818A",
x"B09E808C",
x"AE5D7F7C",
x"ABF47E60",
x"A9717D37",
x"A6EE7C0C",
x"A4857AE5",
x"A24F79CD",
x"A06078CA",
x"9EC577E0",
x"9D827710",
x"9C91765D",
x"9BE375BD",
x"9B5D752F",
x"9AE974AC",
x"9A69742F",
x"99C873B7",
x"98F67347",
x"97EC72DF",
x"96AF7289",
x"95487245",
x"93CB721C",
x"924A720A",
x"90DF7210",
x"8F987226",
x"8E867245",
x"8DAC7261",
x"8D0B726E",
x"8C98725F",
x"8C3E722B",
x"8BDF71C8",
x"8B5D712D",
x"8A917052",
x"89566F31",
x"878A6DC7",
x"85156C10",
x"81E96A0D",
x"7E0767C5",
x"7983653F",
x"747F628D",
x"6F2E5FC5",
x"69D15D01",
x"64AB5A5F",
x"600357FB",
x"5C1355F0",
x"590D5451",
x"570C532C",
x"56175281",
x"56225247",
x"5709526D",
x"589F52DE",
x"5AAA537F",
x"5CF1543A",
x"5F3B54FD",
x"615E55B6",
x"63385663",
x"64B85701",
x"65D95797",
x"66A45828",
x"672758BD",
x"6778595A",
x"67B059FE",
x"67E25AA5",
x"68245B4C",
x"68805BE7",
x"68FF5C74",
x"69A05CEC",
x"6A5F5D4F",
x"6B345D9E",
x"6C135DE0",
x"6CEE5E1C",
x"6DB55E57",
x"6E5C5E95",
x"6ED25ED7",
x"6F115F18",
x"6F145F52",
x"6ED95F76",
x"6E665F7C",
x"6DC75F59",
x"6D0A5F0A",
x"6C425E8D",
x"6B845DEC",
x"6AE25D35",
x"6A6C5C78",
x"6A2E5BCF",
x"6A2B5B4B",
x"6A655AFD",
x"6ACF5AF1",
x"6B615B2C",
x"6C075BA8",
x"6CB45C59",
x"6D545D2E",
x"6DDE5E0E",
x"6E4A5EE4",
x"6E945F9D",
x"6EC56028",
x"6EE3607A",
x"6EF96095",
x"6F14607D",
x"6F41603F",
x"6F895FE9",
x"6FEF5F90",
x"70775F45",
x"71205F15",
x"71DF5F0B",
x"72AE5F2B",
x"73805F70",
x"74495FD2",
x"75006043",
x"759760B5",
x"76096118",
x"764C6163",
x"7660618D",
x"76466194",
x"7601617E",
x"759A6156",
x"751D6128",
x"74966101",
x"741460F2",
x"73A56100",
x"73586134",
x"7330618A",
x"733261FE",
x"735E6283",
x"73A7630A",
x"74046387",
x"746663EA",
x"74BD642B",
x"74F96441",
x"7513642B",
x"750263EC",
x"74C86389",
x"7468630A",
x"73EC627C",
x"736061E9",
x"72CF615F",
x"724460E6",
x"71C56088",
x"715B604D",
x"71036039",
x"70BC604D",
x"70836087",
x"705160DF",
x"7021614C",
x"6FF061C2",
x"6FBB6231",
x"6F80628A",
x"6F4262C1",
x"6F0662CB",
x"6ECE62A1",
x"6E9E6245",
x"6E7C61BB",
x"6E63610D",
x"6E56604B",
x"6E4E5F81",
x"6E445EC2",
x"6E2E5E15",
x"6E035D83",
x"6DB45D0E",
x"6D375CB2",
x"6C835C66",
x"6B905C1E",
x"6A5B5BCD",
x"68E55B66",
x"67315ADD",
x"65495A2E",
x"633B5953",
x"6114584F",
x"5EE65726",
x"5CC555E6",
x"5AC25498",
x"58F0534A",
x"575B520C",
x"561050ED",
x"55174FFB",
x"54734F43",
x"54234ED0",
x"54234EAA",
x"54694ED6",
x"54EE4F51",
x"55A35018",
x"567C511D",
x"576C5251",
x"5865539F",
x"595F54F0",
x"5A51562C",
x"5B345740",
x"5C06581B",
x"5CC758B2",
x"5D795907",
x"5E205921",
x"5EBF590B",
x"5F5E58DA",
x"5FFF58A4",
x"60A6587A",
x"6155586B",
x"62105884",
x"62D458C5",
x"639E5928",
x"646D59A2",
x"653D5A24",
x"66065A9C",
x"66C45B00",
x"67705B42",
x"68065B60",
x"68805B5C",
x"68D65B3D",
x"69095B12",
x"69135AE4",
x"68F75AC3",
x"68B75AB9",
x"68595ACC",
x"67E85AFA",
x"676E5B43",
x"66F95B9F",
x"66995C04",
x"66595C67",
x"664A5CC3",
x"66705D14",
x"66D45D55",
x"67735D8A",
x"684A5DB8",
x"694C5DE6",
x"6A6F5E18",
x"6BA05E56",
x"6CD15EA4",
x"6DF25F00",
x"6EFA5F69",
x"6FE05FDD",
x"70A66056",
x"714960CE",
x"71D5613E",
x"724E61A1",
x"72BF61F6",
x"732D6239",
x"739A626A",
x"7403628B",
x"7465629B",
x"74B5629E",
x"74EA6297",
x"74FA6289",
x"74E06277",
x"749A6266",
x"742E6259",
x"73A76252",
x"73116253",
x"7282625C",
x"7207626A",
x"71B06279",
x"71836281",
x"7183627E",
x"71AA6268",
x"71EB6237",
x"723761E8",
x"727C617A",
x"72AB60F3",
x"72B76059",
x"72975FB7",
x"724C5F1A",
x"71D95E90",
x"71455E25",
x"709B5DE3",
x"6FE95DD0",
x"6F375DEC",
x"6E8F5E32",
x"6DF65E9A",
x"6D735F14",
x"6D075F94",
x"6CB56007",
x"6C806063",
x"6C69609B",
x"6C7360AB",
x"6CA06091",
x"6CEE6052",
x"6D585FF7",
x"6DDC5F8D",
x"6E6C5F21",
x"6EFC5EC1",
x"6F7C5E77",
x"6FDC5E4C",
x"700D5E42",
x"70075E59",
x"6FC25E8A",
x"6F3F5ECB",
x"6E835F0E",
x"6D9B5F48",
x"6C945F69",
x"6B7D5F67",
x"6A665F3E",
x"69595EE9",
x"685F5E6C",
x"677A5DCC",
x"66A95D15",
x"65E65C53",
x"652B5B94",
x"64725AE3",
x"63B15A49",
x"62EB59CC",
x"6220596B",
x"61555925",
x"609758F4",
x"5FF258D0",
x"5F7558B2",
x"5F2D5894",
x"5F2A5874",
x"5F765857",
x"601A5843",
x"611B5846",
x"627D586D",
x"643D58CA",
x"6654596D",
x"68BA5A5C",
x"6B635B9E",
x"6E3F5D2F",
x"713C5F06",
x"7447610E",
x"774C6335",
x"7A3B6560",
x"7D07677A",
x"7FA8696D",
x"821B6B2B",
x"84626CA8",
x"86866DE3",
x"888B6EDC",
x"8A7C6F9C",
x"8C597026",
x"8E227083",
x"8FCD70BD",
x"914F70DB",
x"929370E1",
x"938A70DA",
x"942A70CA",
x"946970BE",
x"945070C1",
x"93EF70E1",
x"935C7129",
x"92BB71A3",
x"922C7254",
x"91D0733B",
x"91BC744E",
x"91FE757C",
x"929476AD",
x"937077C7",
x"947B78B0",
x"959B7954",
x"96B279A6",
x"97A879A3",
x"986D7956",
x"98FB78CE",
x"9959782C",
x"998F7788",
x"99AF7701",
x"99C976AA",
x"99EA7690",
x"9A1876B1",
x"9A567702",
x"9A9B776B",
x"9ADF77D4",
x"9B127822",
x"9B2C783D",
x"9B227816",
x"9AF077A9",
x"9A9576FE",
x"9A187623",
x"99817531",
x"98DA7440",
x"982E736A",
x"978872C3",
x"96F47257",
x"967D722B",
x"962B7240",
x"9604728A",
x"96107300",
x"964F7393",
x"96BF7434",
x"975674DA",
x"98047576",
x"98B67602",
x"99537678",
x"99C076D1",
x"99E97708",
x"99BC771B",
x"99357708",
x"985976D1",
x"973B767B",
x"95F4760C",
x"94AB7592",
x"937D7516",
x"928B74A6",
x"91EA744A",
x"91A27408",
x"91B273E1",
x"920A73D0",
x"929473CB",
x"933573C7",
x"93D573B6",
x"945D738D",
x"94C37348",
x"950772EB",
x"952F727B",
x"954C7208",
x"957071A6",
x"95B17166",
x"961F715C",
x"96C67192",
x"97A87209",
x"98C072BE",
x"9A0373A3",
x"9B5D74A1",
x"9CBC75A3",
x"9E0A768D",
x"9F32774E",
x"A02677D7",
x"A0DC781F",
x"A14F782A",
x"A17B7802",
x"A16677B3",
x"A10E774B",
x"A07676DA",
x"9F997665",
x"9E7175F1",
x"9CF17578",
x"9B0574EA",
x"989B7439",
x"95A4734E",
x"9214721A",
x"8DEF7092",
x"89436EB0",
x"84356C7A",
x"7EF96A06",
x"79CE676C",
x"750064CF",
x"70D86253",
x"6D996021",
x"6B755E56",
x"6A875D0D",
x"6AD25C52",
x"6C3A5C28",
x"6E8D5C86",
x"718A5D5C",
x"74E55E90",
x"78556008",
x"7B9A61AD",
x"7E846362",
x"80FC6518",
x"82FA66C4",
x"848D685C",
x"85D269E2",
x"86EA6B57",
x"87F76CBB",
x"89156E10",
x"8A566F58",
x"8BC0708C",
x"8D5071A9",
x"8EFC72A6",
x"90AF737B",
x"925D7423",
x"93F67499",
x"957074DB",
x"96C974EE",
x"97FE74D8",
x"991474A5",
x"9A0B745B",
x"9AE4740C",
x"9B9B73BE",
x"9C2E737E",
x"9C91734E",
x"9CC27334",
x"9CB97331",
x"9C777341",
x"9C017362",
x"9B5F738F",
x"9A9E73C0",
x"99CD73EF",
x"98FE741A",
x"983B743B",
x"9788744E",
x"96EC7452",
x"965F744A",
x"95DD7436",
x"955D741A",
x"94D973FF",
x"944B73EA",
x"93B473DE",
x"931773E1",
x"927B73F1",
x"91EC740B",
x"91707427",
x"9110743D",
x"90CF743E",
x"90AF7425",
x"90AE73E6",
x"90C67383",
x"90F17302",
x"9129726C",
x"916971D2",
x"91AE714A",
x"91F370E5",
x"923970B5",
x"927E70C7",
x"92BE711C",
x"92F671AD",
x"931F7270",
x"93367352",
x"9339743B",
x"93247517",
x"92FA75D4",
x"92C27662",
x"928776BA",
x"925576DB",
x"923876CB",
x"923E7692",
x"926D763C",
x"92CA75D2",
x"93527564",
x"93FE74F9",
x"94C17499",
x"958B744A",
x"964D7410",
x"96F873EB",
x"978073DA",
x"97DA73D8",
x"980873E1",
x"980A73EE",
x"97E773F8",
x"97AB73FB",
x"976273F1",
x"971773DB",
x"96DA73C1",
x"96B373A9",
x"96AB739C",
x"96BF73A5",
x"96EE73CA",
x"972E740B",
x"976E7462",
x"979D74C3",
x"97A47517",
x"97737548",
x"96FB753E",
x"963374EB",
x"951B7443",
x"93BF734E",
x"922F721C",
x"908B70CA",
x"8EF06F7A",
x"8D816E54",
x"8C5A6D75",
x"8B8E6CF3",
x"8B256CD7",
x"8B146D17",
x"8B426D99",
x"8B856E37",
x"8BAB6EC4",
x"8B796F13",
x"8AB96EF9",
x"893F6E5B",
x"86EF6D2A",
x"83C26B6C",
x"7FCF6937",
x"7B4766AB",
x"766A63F9",
x"71916152",
x"6D175EE9",
x"69525CEA",
x"668F5B77",
x"64FF5AA6",
x"64BA5A7B",
x"65B85AF0",
x"67D85BF0",
x"6AE15D5D",
x"6E8A5F15",
x"728C60F7",
x"769D62E2",
x"7A8664BB",
x"7E216676",
x"815D680C",
x"843C6982",
x"86D16AE2",
x"89316C3B",
x"8B796D9D",
x"8DBE6F14",
x"900D70A6",
x"9266724E",
x"94C27406",
x"971075BC",
x"9939775A",
x"9B2E78D0",
x"9CDD7A06",
x"9E3C7AF4",
x"9F4C7B8F",
x"A0147BD9",
x"A0A27BD9",
x"A1087B9F",
x"A15F7B3C",
x"A1B67AC6",
x"A2257A50",
x"A2B979ED",
x"A37879A8",
x"A4677988",
x"A57B7990",
x"A6A579BA",
x"A7CA79F7",
x"A8C77A34",
x"A9747A61",
x"A9A57A64",
x"A9367A2A",
x"A80879AA",
x"A60F78E0",
x"A35377D0",
x"9FEC768C",
x"9C087530",
x"97EA73DC",
x"93D772B6",
x"901571DA",
x"8CE5715F",
x"8A6D7151",
x"88C671AB",
x"87EC725C",
x"87BF734A",
x"8814744B",
x"88AF753B",
x"895975F9",
x"89DC7668",
x"8A11767B",
x"89E77630",
x"895A7593",
x"887C74B9",
x"876973BD",
x"864572BB",
x"853571CD",
x"84587106",
x"83BF706F",
x"83727009",
x"83696FD1",
x"83916FB7",
x"83CF6FAE",
x"84006FA4",
x"840B6F8F",
x"83D86F65",
x"83606F26",
x"82AD6ED7",
x"81D66E86",
x"81066E48",
x"80726E33",
x"80526E5F",
x"80DF6EE2",
x"82426FCA",
x"8494711D",
x"87D572DA",
x"8BE974EC",
x"909B773C",
x"95A579A3",
x"9AAF7BF8",
x"9F627E0F",
x"A3707FC5",
x"A69980FB",
x"A8B981A2",
x"A9C681B7",
x"A9CF814A",
x"A8FA8070",
x"A7817F49",
x"A5A17DFB",
x"A3987CA3",
x"A1A17B60",
x"9FE17A43",
x"9E787956",
x"9D6D7899",
x"9CBD7806",
x"9C57778F",
x"9C247726",
x"9C0776C0",
x"9BE47657",
x"9BA575E5",
x"9B387571",
x"9A9474FF",
x"99B5749A",
x"98A4744B",
x"976A741A",
x"961A7409",
x"94BF7415",
x"93697431",
x"921B744E",
x"90CE7455",
x"8F74742C",
x"8DF373B9",
x"8C2872E5",
x"89F4719F",
x"87376FDB",
x"83DF6D9D",
x"7FEA6AF5",
x"7B6F67F9",
x"769464D2",
x"719A61AB",
x"6CCF5EB3",
x"68835C1B",
x"65085A0B",
x"629A589F",
x"616557EA",
x"617557E9",
x"62BA588C",
x"650459BB",
x"68145B4C",
x"6B9A5D18",
x"6F475EF7",
x"72D260C8",
x"76076272",
x"78CB63E9",
x"7B16652F",
x"7CFA6655",
x"7EA1676C",
x"8037688E",
x"81ED69D8",
x"83F26B5B",
x"86606D24",
x"894B6F37",
x"8CAB7188",
x"906A7403",
x"9466768B",
x"986D78FE",
x"9C4F7B37",
x"9FDA7D16",
x"A2E47E82",
x"A54D7F68",
x"A7047FCA",
x"A8087FAD",
x"A8647F29",
x"A8367E5B",
x"A7A17D67",
x"A6D07C71",
x"A5F67B9C",
x"A5397B04",
x"A4C07AB6",
x"A4A57ABA",
x"A4F37B08",
x"A5A37B8F",
x"A6A97C39",
x"A7E77CEE",
x"A93B7D96",
x"AA7D7E20",
x"AB8B7E81",
x"AC477EB3",
x"AC9E7EB9",
x"AC877E9B",
x"AC077E61",
x"AB2B7E15",
x"AA0C7DBC",
x"A8C77D59",
x"A77B7CED",
x"A6457C7A",
x"A53C7BFB",
x"A4747B77",
x"A3F47AEF",
x"A3BF7A6F",
x"A3C97A05",
x"A40479BA",
x"A45F799C",
x"A4C079B3",
x"A5177A02",
x"A5547A85",
x"A5717B30",
x"A5717BF8",
x"A55E7CCA",
x"A54D7D95",
x"A5547E4F",
x"A58D7EED",
x"A60B7F6E",
x"A6DC7FD9",
x"A7FE8033",
x"A9668085",
x"AAFA80D9",
x"AC998132",
x"AE1E8191",
x"AF6481F2",
x"B04A824D",
x"B0BF8297",
x"B0BC82C6",
x"B04982D1",
x"AF7A82B6",
x"AE708278",
x"AD4A821B",
x"AC2D81AB",
x"AB318133",
x"AA6780C2",
x"A9D68060",
x"A97B8011",
x"A9477FD6",
x"A9287FA9",
x"A9077F84",
x"A8D17F59",
x"A87A7F20",
x"A7F77ED7",
x"A7497E77",
x"A6777E04",
x"A58A7D87",
x"A48F7D09",
x"A3947C96",
x"A2A17C39",
x"A1BB7BF5",
x"A0E17BCA",
x"A0117BB4",
x"9F407BA9",
x"9E667B99",
x"9D777B78",
x"9C707B39",
x"9B4F7AD7",
x"9A187A50",
x"98D379A8",
x"978A78E8",
x"9646781C",
x"9510774E",
x"93E57683",
x"92BF75BE",
x"918D74F8",
x"903B7423",
x"8EB27331",
x"8CDA7213",
x"8AAA70BB",
x"881B6F27",
x"853F6D5B",
x"82316B68",
x"7F206968",
x"7C42677F",
x"79D665D3",
x"7818648D",
x"773A63CB",
x"775F63A7",
x"7896642D",
x"7ADB655C",
x"7E116728",
x"820E6979",
x"869A6C31",
x"8B736F2A",
x"905C7241",
x"951C7555",
x"998D7848",
x"9D917B05",
x"A1267D7E",
x"A45D7FAD",
x"A7528199",
x"AA30834D",
x"AD2B84D9",
x"B0758650",
x"B43387C8",
x"B87A894D",
x"BD498AEC",
x"C2888CA2",
x"C8068E6C",
x"CD819039",
x"D2AA91F4",
x"D7369384",
x"DADD94D6",
x"DD7195DB",
x"DEDE968A",
x"DF2E96EC",
x"DE8C9710",
x"DD3B9711",
x"DB929711",
x"D9E89730",
x"D8959789",
x"D7DA9831",
x"D7E1992D",
x"D8B79A73",
x"DA4A9BF1",
x"DC6E9D82",
x"DEE49F00",
x"E162A046",
x"E3A3A12D",
x"E569A19F",
x"E686A18C",
x"E6E4A0F6",
x"E6809FEB",
x"E5769E86",
x"E3E99CE8",
x"E20F9B36",
x"E01A9996",
x"DE439829",
x"DCAD9709",
x"DB769647",
x"DAA695E5",
x"DA3495E2",
x"DA0B962D",
x"DA0896B3",
x"DA05975C",
x"D9DD9810",
x"D97498B8",
x"D8B79940",
x"D7A4999C",
x"D64799C4",
x"D4B699BB",
x"D30F9985",
x"D172992A",
x"CFFF98B8",
x"CECB983A",
x"CDE297BA",
x"CD469741",
x"CCEA96CF",
x"CCBC9669",
x"CCA7960C",
x"CC9595B3",
x"CC749559",
x"CC3994FC",
x"CBE19497",
x"CB6F942E",
x"CAEB93BE",
x"CA5E934B",
x"C9D392D8",
x"C94C9266",
x"C8C691F2",
x"C837917A",
x"C79690F6",
x"C6D0905F",
x"C5D68FAA",
x"C49E8ED2",
x"C3288DD5",
x"C17A8CB8",
x"BFAB8B84",
x"BDD18A4F",
x"BC0F8931",
x"BA888842",
x"B95A87A1",
x"B899875E",
x"B854878A",
x"B88A8822",
x"B92D891D",
x"BA298A63",
x"BB638BD6",
x"BCBD8D55",
x"BE1F8EBE",
x"BF788FF6",
x"C0C090EC",
x"C1F7919A",
x"C3239209",
x"C4549247",
x"C599926C",
x"C6FF9293",
x"C88F92D1",
x"CA499334",
x"CC2593C7",
x"CE159480",
x"CFFC9554",
x"D1B79629",
x"D31C96DE",
x"D3F89751",
x"D412975E",
x"D33496E0",
x"D12A95BD",
x"CDC693DC",
x"C8EB9134",
x"C2928DC2",
x"BACC8997",
x"B1C984C9",
x"A7D97F84",
x"9D6279FC",
x"92DD746B",
x"88D26F16",
x"7FBC6A38",
x"780C660E",
x"721162C2",
x"6DF9606E",
x"6BC55F18",
x"6B555EB1",
x"6C685F18",
x"6EA36022",
x"71A76198",
x"75176349",
x"78A46509",
x"7C1666B5",
x"7F4B683E",
x"823C69A4",
x"84F96AF3",
x"879A6C3F",
x"8A386DA1",
x"8CF06F2B",
x"8FCF70EB",
x"92D572E1",
x"95F474FF",
x"99187731",
x"9C217958",
x"9EF07B51",
x"A16A7D02",
x"A37D7E51",
x"A5217F36",
x"A65A7FB2",
x"A7337FD0",
x"A7BF7FA6",
x"A8117F4D",
x"A83C7EE0",
x"A84C7E6E",
x"A84C7E09",
x"A83A7DB9",
x"A8197D78",
x"A7E37D46",
x"A7957D19",
x"A72F7CED",
x"A6B57CBF",
x"A6307C91",
x"A5AC7C6B",
x"A5357C57",
x"A4D67C5D",
x"A4987C81",
x"A4807CC7",
x"A4887D29",
x"A4AC7D9E",
x"A4E47E14",
x"A5237E7E",
x"A5607ECF",
x"A5927EF8",
x"A5B87EFA",
x"A5CD7ED6",
x"A5D47E94",
x"A5CF7E3F",
x"A5B97DE3",
x"A58F7D88",
x"A54D7D30",
x"A4E77CDB",
x"A4527C81",
x"A3827C16",
x"A2747B8E",
x"A1267AE1",
x"9FA47A0C",
x"9DFB7915",
x"9C467808",
x"9AA176F9",
x"992C7601",
x"98037539",
x"973B74B4",
x"96E27483",
x"96FB74AC",
x"9781752A",
x"986475EE",
x"998E76E2",
x"9AE777EC",
x"9C5578F1",
x"9DC079D7",
x"9F157A89",
x"A0437AFC",
x"A13F7B2C",
x"A1FE7B1B",
x"A27A7AD3",
x"A2AE7A63",
x"A29479D8",
x"A2297943",
x"A16E78B0",
x"A0647826",
x"9F1777A9",
x"9D907736",
x"9BE776CA",
x"9A32765E",
x"988E75EA",
x"97157565",
x"95E274D0",
x"95067426",
x"948D7371",
x"947A72B6",
x"94C97202",
x"956D7164",
x"965270E9",
x"9760709F",
x"987D708A",
x"999170B0",
x"9A81710D",
x"9B3C7196",
x"9BAE723D",
x"9BCD72EE",
x"9B927395",
x"9AFE741F",
x"9A17747B",
x"98E974A0",
x"97857488",
x"96047434",
x"947A73AD",
x"92F972FE",
x"918E7233",
x"903F7157",
x"8F067073",
x"8DCF6F8C",
x"8C816E9E",
x"8AFD6DA4",
x"89226C93",
x"86D86B61",
x"84136A03",
x"80D66879",
x"7D3C66C5",
x"797064F6",
x"75AD631E",
x"7231615C",
x"6F445FCB",
x"6D1D5E8A",
x"6BE65DB3",
x"6BB45D56",
x"6C835D7A",
x"6E345E18",
x"709A5F22",
x"7378607E",
x"768F6211",
x"79A263B9",
x"7C866560",
x"7F1866EC",
x"814F684F",
x"832D6984",
x"84C46A8A",
x"862E6B6B",
x"87866C2E",
x"88E36CE1",
x"8A586D8D",
x"8BE96E3E",
x"8D986EF9",
x"8F5A6FC4",
x"912470A0",
x"92E9718D",
x"949C728A",
x"96367390",
x"97B37497",
x"990F7597",
x"9A4C7682",
x"9B66774A",
x"9C5977E4",
x"9D217844",
x"9DB57864",
x"9E0D7841",
x"9E2277E5",
x"9DF0775B",
x"9D7876B6",
x"9CC5760C",
x"9BE07572",
x"9ADC74FE",
x"99CC74B9",
x"98C274A9",
x"97CD74CA",
x"96FB7510",
x"9653756B",
x"95DA75C7",
x"95947616",
x"9581764A",
x"95A57661",
x"96037662",
x"96A17658",
x"97847657",
x"98AF7671",
x"9A2176B6",
x"9BD37731",
x"9DB577E4",
x"9FB178C7",
x"A1AB79C7",
x"A3847AD0",
x"A51C7BC4",
x"A6577C8E",
x"A71E7D16",
x"A7637D51",
x"A7247D3A",
x"A6667CD7",
x"A5397C32",
x"A3B37B5D",
x"A1EB7A6B",
x"A0007971",
x"9E0A787E",
x"9C24779C",
x"9A6476D2",
x"98DF7623",
x"97A2758B",
x"96B87508",
x"96247492",
x"95E67426",
x"95F673C3",
x"96457368",
x"96C17315",
x"975572D0",
x"97E7729C",
x"9867727F",
x"98C2727C",
x"98EE7297",
x"98E972D1",
x"98B47325",
x"9858738C",
x"97E273FF",
x"975C7472",
x"96D274D8",
x"96497526",
x"95C27551",
x"953E7552",
x"94B87527",
x"942F74D4",
x"93A7745E",
x"932273D2",
x"92B17341",
x"926272B9",
x"92457247",
x"926A71F8",
x"92DA71CF",
x"939571D1",
x"948D71F6",
x"95AB7237",
x"96CF7286",
x"97D872D8",
x"98A17321",
x"990E735C",
x"990F7380",
x"989E7392",
x"97C5738F",
x"9697737E",
x"952F7362",
x"93AC733E",
x"92297313",
x"90B572DC",
x"8F567295",
x"8E087233",
x"8CBC71AA",
x"8B5C70F4",
x"89CC7003",
x"87FD6ED8",
x"85DF6D6F",
x"83726BD1",
x"80C36A09",
x"7DF06828",
x"7B1D6649",
x"78766487",
x"762B62FD",
x"746561C9",
x"734B6104",
x"72F260BF",
x"73656106",
x"74A361D9",
x"7699632E",
x"792E64F3",
x"7C42670A",
x"7FAF6954",
x"83536BAE",
x"870D6DFA",
x"8AC5701D",
x"8E667208",
x"91E473B0",
x"953B751C",
x"98647655",
x"9B63776F",
x"9E39787C",
x"A0EA7992",
x"A37A7ABC",
x"A5EA7C01",
x"A83F7D63",
x"AA777ED6",
x"AC978049",
x"AE9581AC",
x"B07582E8",
x"B22883EA",
x"B3A384A2",
x"B4D68505",
x"B5AF8512",
x"B61C84CF",
x"B6128443",
x"B58B8380",
x"B4888295",
x"B3178199",
x"B14A809B",
x"AF427FAB",
x"AD1B7ED4",
x"AAFA7E1E",
x"A8F77D8B",
x"A7267D1C",
x"A5947CCD",
x"A4407C98",
x"A3267C77",
x"A23C7C63",
x"A1737C5A",
x"A0C67C5B",
x"A0337C67",
x"9FBF7C82",
x"9F767CB2",
x"9F637CF8",
x"9F947D5B",
x"A0117DDA",
x"A0D67E6E",
x"A1D67F0B",
x"A2FA7FA8",
x"A41F8030",
x"A5228092",
x"A5DD80BC",
x"A63580A2",
x"A618803F",
x"A5857F95",
x"A4917EB2",
x"A3597DA6",
x"A20A7C91",
x"A0DA7B8E",
x"9FFA7ABC",
x"9F957A36",
x"9FCF7A12",
x"A0B07A58",
x"A2397B09",
x"A44D7C16",
x"A6C67D67",
x"A96E7EDE",
x"AC0E8056",
x"AE6981AF",
x"B05382C9",
x"B1A6838B",
x"B24F83EC",
x"B24783E6",
x"B19E8381",
x"B06D82CD",
x"AED981DD",
x"AD0A80CC",
x"AB257FAC",
x"A94D7E96",
x"A79F7D98",
x"A62B7CC0",
x"A4FA7C16",
x"A4127BA2",
x"A3717B67",
x"A3157B63",
x"A2FA7B95",
x"A31C7BFB",
x"A37B7C8C",
x"A40F7D3F",
x"A4D47E05",
x"A5BF7ECD",
x"A6BD7F88",
x"A7BD8025",
x"A8A88096",
x"A96480D0",
x"A9DC80CF",
x"AA018094",
x"A9CC8023",
x"A93C7F8A",
x"A85D7ED6",
x"A73F7E12",
x"A5FD7D4D",
x"A4AB7C94",
x"A3617BEB",
x"A2307B5B",
x"A11F7AE1",
x"A02B7A79",
x"9F487A1F",
x"9E5D79C6",
x"9D4D795E",
x"9BF678D4",
x"9A347815",
x"97E77706",
x"94F97597",
x"915D73B4",
x"8D157157",
x"88326E80",
x"82D96B42",
x"7D3867BB",
x"77906415",
x"72266087",
x"6D425D48",
x"69275A8E",
x"660C5888",
x"64195757",
x"63615705",
x"63DE578F",
x"657558DC",
x"67F95AC3",
x"6B2E5D12",
x"6ED55F98",
x"72A8621F",
x"76706484",
x"79FD66A7",
x"7D35687A",
x"800969FD",
x"827E6B3B",
x"84A76C45",
x"869D6D31",
x"887D6E14",
x"8A636F00",
x"8C677002",
x"8E9A711F",
x"91007255",
x"939A73A5",
x"965F7505",
x"9943766C",
x"9C3877D4",
x"9F317933",
x"A21C7A85",
x"A4F07BC4",
x"A7A27CEF",
x"AA287E05",
x"AC7A7F04",
x"AE8E7FEE",
x"B06180C5",
x"B1EB8188",
x"B32B8239",
x"B41E82D9",
x"B4CA8367",
x"B53883E4",
x"B56D8450",
x"B57A84A9",
x"B56B84EE",
x"B54C851E",
x"B5288535",
x"B5028535",
x"B4DE851C",
x"B4B584F0",
x"B48184B2",
x"B43A8467",
x"B3D78412",
x"B35383BB",
x"B2AC8361",
x"B1E78308",
x"B10B82B2",
x"B025825D",
x"AF438207",
x"AE7081AD",
x"ADB2814F",
x"AD1180EA",
x"AC84807E",
x"AC04800E",
x"AB827F99",
x"AAF67F25",
x"AA507EB5",
x"A9917E4C",
x"A8C07DEE",
x"A7EB7D9F",
x"A7307D63",
x"A6AB7D3C",
x"A67B7D2D",
x"A6B97D37",
x"A7747D5B",
x"A8AB7D95",
x"AA477DE3",
x"AC297E3D",
x"AE1F7EA0",
x"AFFB7F04",
x"B18A7F63",
x"B2A27FB6",
x"B3307FFE",
x"B32F8039",
x"B2B28068",
x"B1D68092",
x"B0CC80B9",
x"AFBF80E1",
x"AEDC810C",
x"AE3D8139",
x"ADF78160",
x"AE01817A",
x"AE47817A",
x"AEAE8154",
x"AF0B8100",
x"AF3D8075",
x"AF287FB6",
x"AEBC7EC9",
x"ADFB7DBC",
x"ACF57CA2",
x"ABC77B95",
x"AA997AAF",
x"A9957A08",
x"A8E679B4",
x"A8A979C3",
x"A8F87A36",
x"A9DA7B09",
x"AB4A7C33",
x"AD327DA0",
x"AF7B7F39",
x"B20480E7",
x"B4A68295",
x"B747842F",
x"B9CA85A9",
x"BC2086FD",
x"BE408828",
x"C023892C",
x"C1CC8A10",
x"C3328AD2",
x"C44E8B74",
x"C50C8BEF",
x"C54E8C32",
x"C4EB8C2A",
x"C3B68BB9",
x"C17F8AC5",
x"BE1C8932",
x"B97286EC",
x"B37E83E7",
x"AC54802C",
x"A4247BD1",
x"9B3C76F8",
x"91FB71D8",
x"88D56CB1",
x"803967C5",
x"78966358",
x"72445FA2",
x"6D865CD2",
x"6A7F5AFE",
x"69315A33",
x"69835A61",
x"6B425B70",
x"6E2D5D33",
x"71F65F7E",
x"7654621F",
x"7AFE64E5",
x"7FBF67A7",
x"84666A48",
x"88D66CB4",
x"8CFE6EE2",
x"90D870D2",
x"945F7290",
x"979A7426",
x"9A8B75A3",
x"9D387716",
x"9FA27889",
x"A1CD7A03",
x"A3BB7B81",
x"A56A7CFA",
x"A6E07E63",
x"A81E7FAC",
x"A92B80C6",
x"AA0B81A1",
x"AAC78233",
x"AB67827A",
x"ABF7827A",
x"AC7D823F",
x"AD0281DA",
x"AD8F8161",
x"AE2F80EB",
x"AEE1808E",
x"AFA98059",
x"B0858051",
x"B16D807B",
x"B25380CF",
x"B32B813C",
x"B3E081B5",
x"B4608226",
x"B49C8282",
x"B48882BF",
x"B41E82D6",
x"B36382C9",
x"B26182A1",
x"B12C8267",
x"AFDD8228",
x"AE9281F1",
x"AD6481CC",
x"AC6E81C0",
x"ABBF81D0",
x"AB5E81FB",
x"AB4C823D",
x"AB7E828E",
x"ABE182E6",
x"AC608338",
x"ACDD837A",
x"AD4283A5",
x"AD7A83AC",
x"AD74838C",
x"AD29833F",
x"AC9882C2",
x"ABC68215",
x"AAC0813F",
x"A9968049",
x"A85C7F3F",
x"A7257E32",
x"A6047D33",
x"A50B7C56",
x"A44C7BAF",
x"A3CD7B49",
x"A3957B30",
x"A3A47B64",
x"A3EE7BDB",
x"A46A7C86",
x"A4FE7D4D",
x"A5927E11",
x"A60A7EAF",
x"A6497F0B",
x"A63C7F0F",
x"A5D27EAD",
x"A5057DE4",
x"A3DD7CC1",
x"A2697B60",
x"A0C579E1",
x"9F0E786F",
x"9D667731",
x"9BE67647",
x"9AA675C4",
x"99B275B0",
x"990875FF",
x"98A27699",
x"9871775B",
x"98667822",
x"987178C6",
x"988D792A",
x"98B27941",
x"98E77909",
x"9938788D",
x"99AE77E7",
x"9A527734",
x"9B297696",
x"9C2E7626",
x"9D5275F5",
x"9E81760B",
x"9FA27660",
x"A09A76E2",
x"A155777C",
x"A1C37818",
x"A1E478A0",
x"A1BF7909",
x"A164794D",
x"A0EB7972",
x"A0667983",
x"9FE4798E",
x"9F67799B",
x"9EE379AD",
x"9E3F79C0",
x"9D5679C1",
x"9BFD799B",
x"9A0B792C",
x"9764785B",
x"93FB7713",
x"8FDA754A",
x"8B287306",
x"86217061",
x"81136D82",
x"7C596A9A",
x"784E67E2",
x"753F6590",
x"736663D2",
x"72DF62C5",
x"73AA6277",
x"75A762E2",
x"789A63ED",
x"7C396577",
x"80316752",
x"842E694F",
x"87ED6B44",
x"8B386D10",
x"8DF66E9A",
x"901D6FD8",
x"91B970CE",
x"92EA7185",
x"93D0720F",
x"9492727F",
x"955272E8",
x"9628735B",
x"972273E2",
x"98457480",
x"998B7536",
x"9AEA75FC",
x"9C5076CA",
x"9DAE7796",
x"9EF37857",
x"A0127902",
x"A1057996",
x"A1C37A0C",
x"A24C7A65",
x"A29C7AA5",
x"A2B87AC9",
x"A29E7AD7",
x"A2557ACD",
x"A1E37AAF",
x"A14D7A79",
x"A09F7A2D",
x"9FE479C9",
x"9F27794E",
x"9E7478BD",
x"9DD7781B",
x"9D5A776B",
x"9D0176B7",
x"9CD07606",
x"9CC37561",
x"9CD574CE",
x"9CFA7455",
x"9D2973F9",
x"9D5673BB",
x"9D74739A",
x"9D767395",
x"9D5673A6",
x"9D0D73C6",
x"9C9773EE",
x"9BF47415",
x"9B257431",
x"9A2F743D",
x"9918742F",
x"97E97402",
x"96A873B6",
x"9562734B",
x"942172CA",
x"92F1723B",
x"91DD71AB",
x"90ED7129",
x"902570C1",
x"8F87707E",
x"8F117062",
x"8EBB7070",
x"8E7E70A1",
x"8E5270E8",
x"8E2A7134",
x"8DFE7178",
x"8DCB71A1",
x"8D8D71A6",
x"8D467183",
x"8CFD7139",
x"8CB470D1",
x"8C73705A",
x"8C3E6FE1",
x"8C146F79",
x"8BF76F30",
x"8BE26F0D",
x"8BCE6F13",
x"8BB46F3E",
x"8B8A6F86",
x"8B4C6FDC",
x"8AF67034",
x"8A86707F",
x"89FC70AE",
x"896070BB",
x"88BB70A3",
x"88177065",
x"87807008",
x"87036F94",
x"86AE6F16",
x"868B6E99",
x"86A06E29",
x"86F36DCF",
x"87806D93",
x"88426D78",
x"892B6D7C",
x"8A296D9A",
x"8B276DC8",
x"8C0B6DFA",
x"8CBE6E23",
x"8D2A6E38",
x"8D3F6E2E",
x"8CFA6E06",
x"8C5C6DBE",
x"8B6F6D62",
x"8A486CFF",
x"88FC6CA3",
x"87A26C5C",
x"864C6C35",
x"85016C31",
x"83C16C45",
x"827C6C5E",
x"811B6C61",
x"7F816C2A",
x"7D916B97",
x"7B346A8D",
x"785D68FA",
x"751766DE",
x"717C644B",
x"6DBB6168",
x"6A0F5E67",
x"66BF5B88",
x"640D590C",
x"62365730",
x"6161561E",
x"61A155F3",
x"62F256AF",
x"65385840",
x"68475A81",
x"6BE85D3D",
x"6FE2603C",
x"74006344",
x"78186624",
x"7C0E68BB",
x"7FD36AF7",
x"83626CD5",
x"86C16E5F",
x"89F96FA9",
x"8D1470C8",
x"901A71D4",
x"930B72DE",
x"95EA73F1",
x"98B2750F",
x"9B5F7634",
x"9DED775A",
x"A05A7874",
x"A2A67979",
x"A4CF7A63",
x"A6D27B2C",
x"A8AB7BD6",
x"AA517C63",
x"ABBC7CD6",
x"ACDE7D35",
x"ADAB7D82",
x"AE1C7DC1",
x"AE307DF4",
x"ADED7E19",
x"AD5E7E32",
x"AC9C7E3D",
x"ABBD7E3C",
x"AADE7E30",
x"AA197E1E",
x"A9827E09",
x"A9257DF4",
x"A9057DE3",
x"A91E7DD6",
x"A9637DD0",
x"A9C27DD0",
x"AA2B7DD6",
x"AA8C7DE1",
x"AAD97DF4",
x"AB0A7E0C",
x"AB1E7E2C",
x"AB177E56",
x"AAFD7E8A",
x"AAD77EC7",
x"AAAE7F0B",
x"AA847F53",
x"AA5C7F98",
x"AA327FD1",
x"AA047FF8",
x"A9C98004",
x"A97E7FEE",
x"A91E7FB5",
x"A8AB7F57",
x"A8297EDB",
x"A7A47E4C",
x"A7267DB5",
x"A6C57D26",
x"A68A7CB4",
x"A6857C6F",
x"A6BD7C61",
x"A7327C94",
x"A7DF7D05",
x"A8B57DB2",
x"A9A17E8A",
x"AA8B7F7B",
x"AB5E8074",
x"AC08815B",
x"AC778221",
x"ACA582B8",
x"AC918317",
x"AC458342",
x"ABCC833F",
x"AB3B8319",
x"AAA182DE",
x"AA0F8299",
x"A9948254",
x"A933820F",
x"A8EB81C7",
x"A8B68171",
x"A8848101",
x"A8458068",
x"A7E77F9E",
x"A75A7E99",
x"A6957D5E",
x"A5927BF7",
x"A4547A74",
x"A2EA78ED",
x"A167777E",
x"9FE1763E",
x"9E777546",
x"9D4274A5",
x"9C577461",
x"9BC87479",
x"9B9A74E8",
x"9BC9759A",
x"9C48767C",
x"9D007778",
x"9DD57874",
x"9EAB795B",
x"9F677A20",
x"9FF37AB6",
x"A0437B18",
x"A0567B44",
x"A0317B46",
x"9FE17B23",
x"9F777AE8",
x"9F017AA2",
x"9E887A57",
x"9E0A7A0B",
x"9D7A79BA",
x"9CBD795A",
x"9BB378DA",
x"9A357823",
x"98217723",
x"955C75C4",
x"91DA73FB",
x"8DA871C5",
x"88E36F31",
x"83BF6C57",
x"7E836958",
x"797C6665",
x"74FA63AF",
x"71486166",
x"6EA05FB2",
x"6D275EAF",
x"6CEE5E6A",
x"6DE65EDF",
x"6FF35FF7",
x"72E56195",
x"7680638D",
x"7A8665B1",
x"7EBC67DB",
x"82F269E5",
x"87006BBA",
x"8AD06D51",
x"8E566EAD",
x"91976FDC",
x"949C70F6",
x"977A7212",
x"9A437347",
x"9D0874AA",
x"9FDA7646",
x"A2BF7819",
x"A5B57A1D",
x"A8B67C41",
x"ABB37E6D",
x"AE978082",
x"B14F826D",
x"B3C68412",
x"B5E98563",
x"B7AB8659",
x"B90886F1",
x"BA018739",
x"BA9B873F",
x"BAE18717",
x"BADE86D4",
x"BA9F868A",
x"BA2C8643",
x"B9898607",
x"B8B985D3",
x"B7BC85A1",
x"B6918566",
x"B53A8512",
x"B3C0849F",
x"B2358407",
x"B0AB834F",
x"AF3F8281",
x"AE1181B2",
x"AD3F80F8",
x"ACE3806E",
x"AD088028",
x"ADB38036",
x"AEDC809B",
x"B067814F",
x"B2308240",
x"B40C8350",
x"B5CC8460",
x"B73F854D",
x"B84385FD",
x"B8BC8659",
x"B89F865C",
x"B7EE8608",
x"B6BC856E",
x"B52B84A7",
x"B36383CF",
x"B1948305",
x"AFF08264",
x"AEA48200",
x"ADD481E1",
x"AD9C820F",
x"AE078285",
x"AF148336",
x"B0B58417",
x"B2CD8517",
x"B53D862B",
x"B7DE8742",
x"BA898854",
x"BD188958",
x"BF6E8A40",
x"C1748B0A",
x"C31B8BAB",
x"C45D8C1D",
x"C5398C58",
x"C5B68C5A",
x"C5DD8C27",
x"C5BA8BBF",
x"C5598B2E",
x"C4C18A83",
x"C40189CA",
x"C31C8915",
x"C2168873",
x"C0F587EA",
x"BFB68781",
x"BE598735",
x"BCDB8700",
x"BB4286D9",
x"B98F86B3",
x"B7CF868A",
x"B6118657",
x"B46A861C",
x"B2F585DE",
x"B1D485AC",
x"B11F858F",
x"B0ED8597",
x"B14785C8",
x"B22D8627",
x"B38B86A9",
x"B53D8746",
x"B71887E7",
x"B8EA8879",
x"BA7F88E9",
x"BBB58928",
x"BC6E8931",
x"BCA38908",
x"BC6188BB",
x"BBBD8859",
x"BAD687F6",
x"B9CC879F",
x"B8B3875E",
x"B794872F",
x"B65E86FD",
x"B4F486AB",
x"B32C8618",
x"B0D6851B",
x"ADC68395",
x"A9E68174",
x"A5327EB5",
x"9FC87B67",
x"99E077B0",
x"93CB73C4",
x"8DE56FE2",
x"888B6C4D",
x"84176941",
x"80C566ED",
x"7EBC6573",
x"7E0064DA",
x"7E79651B",
x"7FF9661B",
x"824167AE",
x"850D69A6",
x"88216BD1",
x"8B4B6E03",
x"8E697016",
x"916D71F2",
x"9456738C",
x"973174E1",
x"9A0D75FE",
x"9CFD76F2",
x"A00A77D5",
x"A33C78BD",
x"A68D79BE",
x"A9F47AED",
x"AD617C50",
x"B0C67DF1",
x"B40F7FC9",
x"B73281D1",
x"BA2283FE",
x"BCDA863B",
x"BF578874",
x"C1988A97",
x"C3988C91",
x"C5508E53",
x"C6BC8FD1",
x"C7D19100",
x"C88791DD",
x"C8D79266",
x"C8C1929E",
x"C84C9289",
x"C7849231",
x"C68191A2",
x"C56190ED",
x"C4479021",
x"C3518F52",
x"C2A08E94",
x"C2478DF6",
x"C24E8D84",
x"C2B08D49",
x"C35B8D42",
x"C4338D6C",
x"C5158DBC",
x"C5E08E24",
x"C67B8E97",
x"C6D78F0B",
x"C6F78F7D",
x"C6EB8FEF",
x"C6D19066",
x"C6D090F3",
x"C70B919E",
x"C7A09274",
x"C8A59376",
x"CA1594A0",
x"CBE395E0",
x"CDEE9727",
x"D0119858",
x"D222995E",
x"D4059A27",
x"D5A99AAE",
x"D70F9AFB",
x"D8469B1F",
x"D96F9B36",
x"DAAC9B5C",
x"DC1C9BB1",
x"DDD59C45",
x"DFDD9D1F",
x"E2229E34",
x"E4869F71",
x"E6DEA0B1",
x"E8FBA1D3",
x"EAB1A2B3",
x"EBE6A33A",
x"EC8CA35F",
x"ECAAA327",
x"EC5AA2A7",
x"EBBDA1FC",
x"EAF6A148",
x"EA27A0B0",
x"E965A048",
x"E8B1A01D",
x"E7FEA02C",
x"E72EA061",
x"E61FA09C",
x"E4A7A0BA",
x"E2A7A093",
x"E00CA00B",
x"DCD29F08",
x"D90B9D82",
x"D4D59B82",
x"D062991D",
x"CBEA9670",
x"C7A693A5",
x"C3C790E5",
x"C0778E52",
x"BDCD8C0D",
x"BBCE8A28",
x"BA6B88A7",
x"B9858783",
x"B8EE86A5",
x"B87285F4",
x"B7DA854F",
x"B6F58494",
x"B5A083AD",
x"B3C9828B",
x"B171812C",
x"AEAC7F9B",
x"ABA27DF1",
x"A8817C49",
x"A57D7AC1",
x"A2C07975",
x"A0697875",
x"9E7E77C1",
x"9CF07748",
x"9B9876F1",
x"9A39768C",
x"989475F1",
x"966474F2",
x"9374736F",
x"8FA5715A",
x"8AF46EB5",
x"85816B9D",
x"7F8C683C",
x"796864CC",
x"7378618B",
x"6E215EB3",
x"69C05C77",
x"66915AF6",
x"64BD5A39",
x"64445A39",
x"65085ADA",
x"66CC5BF4",
x"69485D57",
x"6C265ED9",
x"6F14604D",
x"71D16197",
x"742862A7",
x"76016379",
x"775B6411",
x"78426480",
x"78D864D8",
x"793E652A",
x"79986583",
x"7A0665EC",
x"7A986665",
x"7B5C66EC",
x"7C4C6777",
x"7D5C67FD",
x"7E7A6876",
x"7F9668D6",
x"809E691D",
x"81846944",
x"8245694F",
x"82DF6942",
x"83566920",
x"83B568F0",
x"840768B8",
x"8455687D",
x"84A56845",
x"84FD6817",
x"855C67F9",
x"85C167EF",
x"86256801",
x"86846835",
x"86D6688D",
x"871B690C",
x"875269AE",
x"87806A70",
x"87AC6B48",
x"87DF6C2B",
x"88206D0C",
x"88776DD9",
x"88E76E86",
x"896C6F02",
x"89FD6F44",
x"8A8D6F44",
x"8B0A6F02",
x"8B5F6E7F",
x"8B7D6DC5",
x"8B596CE3",
x"8AEA6BED",
x"8A386AF7",
x"89496A17",
x"882F695F",
x"870168DF",
x"85D0689D",
x"84B16899",
x"83AF68C9",
x"82D0691E",
x"82156984",
x"817669E6",
x"80EC6A2D",
x"806F6A4C",
x"7FFA6A3B",
x"7F9069FD",
x"7F35699D",
x"7EF7692D",
x"7EE568C5",
x"7F0A687C",
x"7F726866",
x"80216891",
x"811068FD",
x"823169A7",
x"836F6A7D",
x"84AF6B68",
x"85D86C4D",
x"86D56D14",
x"87946DAA",
x"88136E02",
x"88536E1A",
x"88636DF9",
x"88556DAB",
x"883B6D47",
x"88286CDF",
x"88276C86",
x"88396C4B",
x"88596C31",
x"88796C38",
x"888A6C57",
x"88776C7D",
x"88346C9E",
x"87B86CA6",
x"87036C89",
x"86206C3D",
x"851B6BBE",
x"840B6B10",
x"83006A3A",
x"820A6945",
x"81326841",
x"8077673A",
x"7FD2663B",
x"7F32654F",
x"7E89647F",
x"7DC463CF",
x"7CD86345",
x"7BC462E2",
x"7A8A62A7",
x"793E6294",
x"77F262A5",
x"76BC62D5",
x"75B46318",
x"74E36363",
x"744C63A5",
x"73E663CC",
x"739763C5",
x"733F637C",
x"72B862E6",
x"71DD61F7",
x"708F60B1",
x"6EBA5F17",
x"6C5B5D3B",
x"697F5B2F",
x"66475911",
x"62DC56FD",
x"5F75550F",
x"5C475363",
x"5986520C",
x"575C5119",
x"55E75091",
x"55315072",
x"553D50B6",
x"55F65153",
x"57445236",
x"5900534E",
x"5B05548C",
x"5D2E55DA",
x"5F5B572B",
x"6172586E",
x"635F5997",
x"651D5A9E",
x"66A95B7D",
x"68065C31",
x"693E5CBC",
x"6A5E5D27",
x"6B6D5D77",
x"6C795DBB",
x"6D865DFA",
x"6E975E42",
x"6FAB5E9A",
x"70BB5F03",
x"71C15F7E",
x"72B16004",
x"7380608B",
x"74236107",
x"7491616C",
x"74C961AF",
x"74CB61CC",
x"749B61C2",
x"74476197",
x"73DE6158",
x"73726113",
x"731460D6",
x"72D360B2",
x"72BD60AF",
x"72D360D2",
x"73146117",
x"73766177",
x"73ED61E6",
x"74696255",
x"74D962B4",
x"753462FA",
x"7572631E",
x"75916323",
x"75996307",
x"759662D8",
x"7594629B",
x"75A1625F",
x"75C86228",
x"760F6200",
x"767261E6",
x"76E961DA",
x"776B61D9",
x"77E361DF",
x"784561E4",
x"788361E9",
x"789361E8",
x"787061E2",
x"782061D8",
x"77A761CE",
x"770E61C3",
x"766361BC",
x"75AD61B8",
x"74F461B4",
x"744161AF",
x"739761A7",
x"72FA6197",
x"726D617E",
x"71F5615C",
x"71916132",
x"714C6106",
x"712860DC",
x"712860BE",
x"714F60B5",
x"719860C6",
x"720260FA",
x"727F6150",
x"730361C9",
x"7384625F",
x"73F46306",
x"744863AE",
x"74786448",
x"747D64C1",
x"745B6507",
x"7413650E",
x"73AB64CE",
x"73306448",
x"72A86381",
x"721D628D",
x"7198617D",
x"7120606C",
x"70B85F73",
x"70635EA4",
x"70215E11",
x"6FF05DBF",
x"6FCC5DAF",
x"6FAE5DD5",
x"6F905E24",
x"6F6C5E87",
x"6F3E5EED",
x"6F005F46",
x"6EB45F87",
x"6E595FA8",
x"6DF65FAC",
x"6D8F5F98",
x"6D2D5F72",
x"6CD85F41",
x"6C965F0E",
x"6C6D5EDC",
x"6C5E5EAE",
x"6C685E81",
x"6C835E53",
x"6CA75E1E",
x"6CC55DDF",
x"6CCC5D92",
x"6CAD5D38",
x"6C595CD0",
x"6BC25C5D",
x"6AE55BE4",
x"69BC5B67",
x"68545AEA",
x"66B55A74",
x"64F85A04",
x"633459A2",
x"6186594F",
x"600C5911",
x"5EE258ED",
x"5E1E58E6",
x"5DD45902",
x"5E095945",
x"5EBE59AF",
x"5FE95A42",
x"617D5AFA",
x"63655BD2",
x"65875CC5",
x"67CF5DCB",
x"6A245EDC",
x"6C735FF3",
x"6EB16108",
x"70D2621A",
x"72D36321",
x"74B56420",
x"767D6514",
x"783165FC",
x"79D666D6",
x"7B7367A3",
x"7D0B685F",
x"7EA2690A",
x"803869A1",
x"81C56A21",
x"83486A8C",
x"84BA6AE2",
x"86116B24",
x"874C6B5B",
x"88666B87",
x"895F6BB4",
x"8A386BE6",
x"8AF96C23",
x"8BA76C70",
x"8C4E6CD1",
x"8CF46D45",
x"8DA46DCB",
x"8E626E5F",
x"8F326EFF",
x"90136FA4",
x"9100704F",
x"91F370FB",
x"92E271A6",
x"93C37254",
x"948E7302",
x"953973B3",
x"95C17465",
x"96227517",
x"966275C6",
x"9687766B",
x"96A17703",
x"96BD7786",
x"96F077F4",
x"974C784A",
x"97E2788B",
x"98BE78BD",
x"99E678EA",
x"9B5A7916",
x"9D0D794E",
x"9EED7995",
x"A0DC79EB",
x"A2BB7A50",
x"A46A7ABA",
x"A5CA7B22",
x"A6C67B79",
x"A7537BBC",
x"A7747BE0",
x"A73A7BE5",
x"A6C27BD1",
x"A6337BAD",
x"A5B67B85",
x"A5737B68",
x"A58A7B63",
x"A60E7B7C",
x"A7017BBA",
x"A8547C18",
x"A9EB7C8E",
x"AB9C7D0F",
x"AD367D8E",
x"AE8C7DF8",
x"AF747E44",
x"AFD07E6A",
x"AF917E65",
x"AEB97E3C",
x"AD5C7DF4",
x"AB997D99",
x"A99B7D36",
x"A78D7CD7",
x"A59E7C82",
x"A3F77C3C",
x"A2B57C04",
x"A1E77BD7",
x"A1957BAF",
x"A1B37B81",
x"A22E7B49",
x"A2EB7AFE",
x"A3CC7AA3",
x"A4B27A39",
x"A58579C7",
x"A633795A",
x"A6B678FF",
x"A70E78C6",
x"A74278B6",
x"A75E78D8",
x"A774792F",
x"A78D79B0",
x"A7AC7A51",
x"A7D07AFF",
x"A7EE7BA3",
x"A7F77C28",
x"A7D77C7A",
x"A77D7C8C",
x"A6DC7C5B",
x"A5F17BE8",
x"A4C37B3E",
x"A35C7A6E",
x"A1D27983",
x"A036788F",
x"9E977798",
x"9CFB769D",
x"9B5A7599",
x"99A17479",
x"97B1732B",
x"956A719F",
x"92AB6FC4",
x"8F606D96",
x"8B846B1E",
x"87276873",
x"826D65B5",
x"7D94630E",
x"78E060AD",
x"74A15EB9",
x"711B5D5C",
x"6E8F5CA7",
x"6D205CA4",
x"6CDF5D4B",
x"6DBF5E84",
x"6FA46031",
x"72586228",
x"75A06444",
x"793C665F",
x"7CF6685E",
x"809B6A2B",
x"840A6BBE",
x"872C6D14",
x"89FE6E33",
x"8C816F23",
x"8EC36FF0",
x"90D370AB",
x"92C57161",
x"94AB721D",
x"969872EE",
x"989773D8",
x"9AB474E8",
x"9CF0761F",
x"9F4D777C",
x"A1C578FB",
x"A44A7A91",
x"A6CC7C2F",
x"A9357DC0",
x"AB717F2F",
x"AD688068",
x"AF0C815B",
x"B04D81FB",
x"B1268245",
x"B198823B",
x"B1A981E8",
x"B16A8163",
x"B0EA80BA",
x"B03D800A",
x"AF747F5E",
x"AE9E7ECC",
x"ADC47E53",
x"ACF17DF7",
x"AC217DB2",
x"AB567D7A",
x"AA917D41",
x"A9CD7D02",
x"A90C7CB3",
x"A84F7C53",
x"A7987BE4",
x"A6EA7B6D",
x"A6497AFB",
x"A5B57A96",
x"A52F7A4D",
x"A4B67A25",
x"A4477A22",
x"A3E17A43",
x"A3807A81",
x"A3227AD0",
x"A2C77B25",
x"A2737B6F",
x"A2267BA3",
x"A1E67BB6",
x"A1B27BA0",
x"A1887B5D",
x"A1647AEF",
x"A1407A5E",
x"A10F79B2",
x"A0C678F2",
x"A05D7830",
x"9FCD7774",
x"9F1576C8",
x"9E3B7636",
x"9D4B75C1",
x"9C56756F",
x"9B73753E",
x"9AB6752D",
x"9A347539",
x"99F7755E",
x"9A0A759A",
x"9A6975E8",
x"9B0B7644",
x"9BE076AD",
x"9CD57720",
x"9DD5779C",
x"9ECC781F",
x"9FA978A7",
x"A0637932",
x"A0F079BD",
x"A14F7A41",
x"A17E7ABC",
x"A1817B23",
x"A15A7B74",
x"A10B7BA8",
x"A09A7BBA",
x"A00A7BAA",
x"9F627B7B",
x"9EA97B2F",
x"9DEE7AD1",
x"9D3F7A6A",
x"9CAB7A08",
x"9C4579B9",
x"9C1C7988",
x"9C3F7982",
x"9CAF79AD",
x"9D707A0C",
x"9E747A9F",
x"9FAC7B5B",
x"A1017C39",
x"A25A7D28",
x"A39C7E16",
x"A4B57EF2",
x"A5917FAD",
x"A62C803C",
x"A6878098",
x"A6A980BD",
x"A6A180AC",
x"A6788068",
x"A6397FF7",
x"A5E17F5A",
x"A5627E94",
x"A4A17D9E",
x"A37B7C6F",
x"A1C37B01",
x"9F527944",
x"9C01772F",
x"97C274BD",
x"929571F2",
x"8C9A6ED8",
x"86046B86",
x"7F21681B",
x"784864BB",
x"71D9618D",
x"6C2B5EB3",
x"678C5C50",
x"64285A76",
x"621C592E",
x"61615878",
x"61D8584A",
x"63525892",
x"65905936",
x"68545A24",
x"6B5E5B43",
x"6E7C5C84",
x"71865DDA",
x"74625F3E",
x"770160AB",
x"7963621D",
x"7B876391",
x"7D766509",
x"7F3B667C",
x"80DD67E9",
x"82686948",
x"83E26A96",
x"85506BCC",
x"86B96CE9",
x"88206DEB",
x"89836ED1",
x"8AE06F9D",
x"8C347052",
x"8D7470F2",
x"8E987182",
x"8F947200",
x"90607272",
x"90F772D7",
x"9156732D",
x"91847374",
x"918873A7",
x"917173C4",
x"914F73C4",
x"913273A5",
x"91257362",
x"913572FC",
x"91607274",
x"91A571CB",
x"91FA710F",
x"92557048",
x"92A86F86",
x"92E66ED8",
x"93076E4D",
x"93086DF0",
x"92ED6DCD",
x"92BE6DE3",
x"92876E33",
x"92566EB4",
x"92396F5B",
x"92397019",
x"925A70E1",
x"929771A0",
x"92E6724D",
x"933672DC",
x"9374734B",
x"938E7395",
x"937173BB",
x"931773C4",
x"927D73B3",
x"91AE738D",
x"90BB735A",
x"8FBC731C",
x"8ED072DA",
x"8E147295",
x"8D9E7252",
x"8D807215",
x"8DBC71E1",
x"8E5071B9",
x"8F29719F",
x"902E7197",
x"914071A1",
x"923E71BD",
x"930871E2",
x"9387720A",
x"93AB7230",
x"93697245",
x"92C67244",
x"91CC7223",
x"908B71DC",
x"8F1A7172",
x"8D9170E8",
x"8C097043",
x"8A956F8F",
x"894C6ED9",
x"88356E2D",
x"875B6D94",
x"86BB6D17",
x"864F6CBB",
x"860D6C7D",
x"85E66C5B",
x"85C86C4B",
x"85A16C44",
x"85656C3D",
x"85046C2B",
x"847A6C09",
x"83CB6BD1",
x"82FA6B83",
x"82186B23",
x"81376AB1",
x"80696A35",
x"7FC269B8",
x"7F52693F",
x"7F2168CE",
x"7F34686B",
x"7F846814",
x"800967CB",
x"80AE678E",
x"81626758",
x"82106725",
x"82A166F0",
x"830666B7",
x"832B6673",
x"83046623",
x"828665C4",
x"81A76552",
x"806264CC",
x"7EB0642D",
x"7C8E6372",
x"7A026297",
x"77106195",
x"73C7606E",
x"703C5F1F",
x"6C8D5DAC",
x"68DB5C1F",
x"654D5A82",
x"620958EA",
x"5F31576A",
x"5CE55619",
x"5B37550C",
x"5A315457",
x"59CF5405",
x"5A06541C",
x"5AC15498",
x"5BE4556D",
x"5D555688",
x"5EF957D1",
x"60BA5932",
x"62865A8E",
x"64525BD2",
x"66165CED",
x"67CE5DD9",
x"69765E91",
x"6B0C5F1B",
x"6C8C5F7E",
x"6DF05FC6",
x"6F315FFD",
x"704B602B",
x"71386058",
x"71F66088",
x"728760BC",
x"72F360F3",
x"7344612B",
x"73846160",
x"73C76190",
x"741461B9",
x"747861DA",
x"74F761F6",
x"7593620E",
x"76466227",
x"770A6243",
x"77D3626A",
x"7897629F",
x"794B62E8",
x"79E66342",
x"7A6063AF",
x"7AB5642D",
x"7AE664B2",
x"7AF2653A",
x"7ADB65B5",
x"7AA8661B",
x"7A5D6663",
x"7A046683",
x"79A4667C",
x"7944664B",
x"78EC65F7",
x"78A7658B",
x"78796513",
x"7865649A",
x"786D642D",
x"788E63D2",
x"78C1638D",
x"78FF6362",
x"793A634C",
x"79686346",
x"797F634B",
x"79766353",
x"794C635A",
x"7901635F",
x"7898635D",
x"781D6355",
x"77976348",
x"77116335",
x"7697631B",
x"763062FD",
x"75E062D6",
x"75AD62AB",
x"7593627C",
x"7590624C",
x"75A16221",
x"75C26201",
x"75F061F4",
x"762761FC",
x"7666621B",
x"76AD6252",
x"76F76297",
x"774862E4",
x"779B632D",
x"77F06363",
x"78426380",
x"7890637C",
x"78D36353",
x"7909630E",
x"792A62B1",
x"79306248",
x"791761E2",
x"78DB6187",
x"78766143",
x"77EC6118",
x"773E610A",
x"76736113",
x"7597612D",
x"74BA6152",
x"73EC617E",
x"734161AB",
x"72C861D9",
x"728E6207",
x"729D6239",
x"72F36270",
x"738762AE",
x"744962F3",
x"7525633B",
x"76016381",
x"76C563C1",
x"775F63F0",
x"77BE640D",
x"77E06411",
x"77C963FF",
x"778663D5",
x"77236398",
x"76B2634E",
x"764562F7",
x"75E0629A",
x"75866235",
x"752A61C8",
x"74BB614C",
x"742460C1",
x"7348601D",
x"72135F5F",
x"70765E84",
x"6E6D5D8E",
x"6C025C82",
x"69485B6A",
x"66635A4D",
x"637C5939",
x"60BE583A",
x"5E54575C",
x"5C6256A5",
x"5B00561F",
x"5A3E55CC",
x"5A1755AC",
x"5A8055BA",
x"5B5E55F1",
x"5C925649",
x"5DF656B9",
x"5F6B5736",
x"60D257B9",
x"6216583D",
x"632758BF",
x"64035939",
x"64AE59AF",
x"65305A1F",
x"65975A8E",
x"65F05AFA",
x"664B5B63",
x"66AE5BC9",
x"67205C29",
x"67A35C81",
x"68345CCC",
x"68CF5D08",
x"696F5D38",
x"6A115D5C",
x"6AB15D7A",
x"6B4E5D97",
x"6BE95DBD",
x"6C865DF4",
x"6D275E41",
x"6DCE5EA8",
x"6E7C5F2B",
x"6F2D5FC9",
x"6FDC607D",
x"70836141",
x"7119620B",
x"719462D5",
x"71F06397",
x"722A6449",
x"724164E6",
x"723B656A",
x"722365D2",
x"72076618",
x"71F6663F",
x"72006645",
x"7230662A",
x"729165F3",
x"732765A3",
x"73EF6544",
x"74E364DE",
x"75FA647D",
x"7724642D",
x"785663FA",
x"798263EF",
x"7A9D6410",
x"7BA06462",
x"7C8A64E0",
x"7D5B6584",
x"7E136641",
x"7EB7670A",
x"7F4867CC",
x"7FC96877",
x"80386900",
x"80936958",
x"80D2697A",
x"80F36968",
x"80EF6924",
x"80C568BB",
x"8074683A",
x"800167B1",
x"7F70672E",
x"7ECB66BE",
x"7E1A6668",
x"7D656630",
x"7CB16611",
x"7C046603",
x"7B6065FA",
x"7AC565E6",
x"7A3165BC",
x"79A56573",
x"79216507",
x"78AD647C",
x"784B63DA",
x"78066335",
x"77E5629D",
x"77F06227",
x"782761E2",
x"788661D8",
x"7904620B",
x"798E6276",
x"7A116309",
x"7A7463AF",
x"7AA56453",
x"7A9364DE",
x"7A37653F",
x"7997656D",
x"78C26568",
x"77D16537",
x"76E064E8",
x"7614648E",
x"7586643F",
x"754E640A",
x"757263FC",
x"75EF6415",
x"76B56453",
x"77A764A8",
x"78A16504",
x"797F6550",
x"7A1E657D",
x"7A65657D",
x"7A476548",
x"79C464E0",
x"78E7644F",
x"77CC63A4",
x"768D62F2",
x"7547624C",
x"741661C3",
x"730A615F",
x"72276121",
x"71686101",
x"70B860F0",
x"700160DC",
x"6F2560AD",
x"6E0D604F",
x"6CA65FB5",
x"6AF05EDD",
x"68F65DCC",
x"66D55C92",
x"64B45B49",
x"62C15A0E",
x"612E5901",
x"6026583C",
x"5FC757D1",
x"601F57CD",
x"612A582B",
x"62D258DF",
x"64F359D3",
x"67605AF1",
x"69E95C1E",
x"6C625D45",
x"6EA85E53",
x"70A75F43",
x"72586014",
x"73C160C9",
x"74F0616F",
x"75FC620B",
x"76F662A8",
x"77ED6348",
x"78E763EC",
x"79E2648E",
x"7AD26528",
x"7BAA65AE",
x"7C596618",
x"7CD46662",
x"7D106689",
x"7D116690",
x"7CE2667F",
x"7C8E665C",
x"7C2B6635",
x"7BCE6613",
x"7B8365FC",
x"7B5865F6",
x"7B516604",
x"7B686621",
x"7B94664B",
x"7BCB667C",
x"7BFD66AA",
x"7C2066CF",
x"7C2B66E6",
x"7C1D66EC",
x"7BF966E0",
x"7BC566C6",
x"7B8D66A3",
x"7B5C667F",
x"7B3B6662",
x"7B356659",
x"7B4E666D",
x"7B8666A7",
x"7BDF6707",
x"7C52678E",
x"7CDA6838",
x"7D7068F7",
x"7E0E69BF",
x"7EAE6A7D",
x"7F4C6B21",
x"7FE26B9C",
x"80706BDE",
x"80F36BE3",
x"81696BAD",
x"81CF6B3F",
x"82256AA6",
x"826869F2",
x"82946934",
x"82AB687F",
x"82AA67E3",
x"8295676C",
x"82736724",
x"824C6710",
x"8228672D",
x"82146779",
x"821B67EC",
x"8246687C",
x"8298691E",
x"831169C7",
x"83A86A65",
x"84526AEF",
x"84FB6B57",
x"85946B93",
x"86096B9E",
x"864E6B76",
x"86586B1E",
x"862A6AA0",
x"85C66A07",
x"853B6968",
x"849A68D2",
x"83F2685B",
x"83566810",
x"82D567FD",
x"82776826",
x"82426887",
x"82356919",
x"824F69CC",
x"828B6A93",
x"82E36B59",
x"83556C10",
x"83DA6CAB",
x"84706D26",
x"85106D79",
x"85B46DAA",
x"86536DBB",
x"86E06DB4",
x"87526D9C",
x"879D6D78",
x"87B56D4E",
x"87966D21",
x"87426CF2",
x"86BF6CC2",
x"861B6C90",
x"85666C5C",
x"84B26C27",
x"84156BEF",
x"839B6BB5",
x"834B6B7C",
x"83286B42",
x"832B6B0A",
x"83456AD2",
x"83636A99",
x"836F6A5C",
x"83526A17",
x"82F769C2",
x"82496959",
x"813B68CF",
x"7FBF681A",
x"7DD06731",
x"7B6F660B",
x"789D64A1",
x"756962F3",
x"71E56106",
x"6E285EE6",
x"6A545CA8",
x"668D5A64",
x"62FB583C",
x"5FC4564D",
x"5D0C54B5",
x"5AEC538C",
x"597652E3",
x"58B052BA",
x"5890530E",
x"590553C9",
x"59F354D0",
x"5B3D5601",
x"5CC1573C",
x"5E66585F",
x"60145950",
x"61BD5A02",
x"63585A73",
x"64E55AA5",
x"66655AAE",
x"67DE5AA5",
x"69515AA4",
x"6ABE5AC6",
x"6C235B1F",
x"6D795BC0",
x"6EB75CA8",
x"6FD25DD2",
x"70C25F2B",
x"7182609B",
x"720D6203",
x"72656344",
x"72916441",
x"729864E8",
x"7284652A",
x"72636509",
x"723B6490",
x"721863D5",
x"720262F3",
x"71F7620E",
x"71FD6143",
x"721160AF",
x"72306064",
x"7255606C",
x"727C60C3",
x"72A1615D",
x"72C46222",
x"72E862F7",
x"731063BF",
x"73446462",
x"738E64C9",
x"73FA64EC",
x"748D64C8",
x"754C6466",
x"763863D9",
x"77496337",
x"78776297",
x"79AF6214",
x"7AE261C2",
x"7BF961AE",
x"7CE661DD",
x"7D9D6253",
x"7E166306",
x"7E5063E6",
x"7E5564E5",
x"7E2A65EF",
x"7DDD66F2",
x"7D7F67DE",
x"7D1A68A8",
x"7CBA694B",
x"7C6969BF",
x"7C2B6A07",
x"7C066A28",
x"7BFF6A27",
x"7C176A0D",
x"7C5369DF",
x"7CB769A6",
x"7D446969",
x"7DF9692B",
x"7ED568F5",
x"7FD168C7",
x"80DD68A7",
x"81EF6896",
x"82EF6899",
x"83CB68B0",
x"846F68DB",
x"84CC691A",
x"84DC6968",
x"849D69BE",
x"84186A16",
x"835D6A63",
x"82846A9D",
x"81A76AB8",
x"80DD6AAE",
x"803C6A79",
x"7FD26A17",
x"7FA4698D",
x"7FAA68E2",
x"7FD8681E",
x"80166751",
x"804B6686",
x"805F65CB",
x"803F652A",
x"7FDD64AA",
x"7F3A644F",
x"7E5B641A",
x"7D506406",
x"7C316410",
x"7B136431",
x"7A0C6460",
x"792A649B",
x"787564D9",
x"77E96514",
x"77816546",
x"772D656D",
x"76D96581",
x"767A657F",
x"7601655F",
x"7568651D",
x"74AD64B5",
x"73D36427",
x"72DE6372",
x"71D36295",
x"70B56198",
x"6F806081",
x"6E2E5F55",
x"6CB55E1B",
x"6B0C5CDA",
x"69285B98",
x"67095A5C",
x"64B55926",
x"623E5800",
x"5FBD56EA",
x"5D5155ED",
x"5B21550F",
x"59515459",
x"580053D1",
x"5745537F",
x"5729536B",
x"57A95393",
x"58B553F5",
x"5A34548C",
x"5C09554D",
x"5E105629",
x"602D5712",
x"624857FD",
x"644E58DD",
x"663D59AC",
x"68115A6B",
x"69D85B1F",
x"6B985BD0",
x"6D635C8A",
x"6F425D57",
x"713A5E45",
x"734C5F58",
x"75736090",
x"77A461E6",
x"79D2634E",
x"7BED64B8",
x"7DE56610",
x"7FAB6744",
x"81396842",
x"828A6901",
x"839A697C",
x"846D69B5",
x"850A69BA",
x"85796997",
x"85C26962",
x"85EF6931",
x"86096916",
x"86186921",
x"8628695B",
x"863C69C7",
x"86606A5F",
x"86986B1C",
x"86EC6BEC",
x"87606CC2",
x"87F96D8F",
x"88B46E45",
x"89936EDF",
x"8A8D6F58",
x"8BA16FB3",
x"8CC26FF5",
x"8DEA7027",
x"8F107054",
x"90287082",
x"912F70B9",
x"921D70FB",
x"92ED7147",
x"939E719A",
x"942E71EC",
x"94977237",
x"94DA7272",
x"94F47299",
x"94E172A7",
x"94A1729F",
x"94327280",
x"93987254",
x"92D87220",
x"91FA71EC",
x"910E71C0",
x"902171A1",
x"8F437193",
x"8E867195",
x"8DF471A0",
x"8D9871B0",
x"8D7471BB",
x"8D8771BE",
x"8DC871B0",
x"8E2A718D",
x"8E9B7158",
x"8F0B7113",
x"8F6A70C3",
x"8FA97070",
x"8FBF7024",
x"8FA76FE4",
x"8F606FB1",
x"8EEF6F92",
x"8E5A6F7F",
x"8DAC6F78",
x"8CED6F73",
x"8C286F69",
x"8B636F55",
x"8AA76F30",
x"89F76EF9",
x"89596EAE",
x"88D26E52",
x"88656DEC",
x"88156D82",
x"87EC6D1C",
x"87EF6CBF",
x"88216C78",
x"88886C4B",
x"89256C3E",
x"89F66C57",
x"8AF06C94",
x"8C076CF5",
x"8D276D73",
x"8E386E03",
x"8F1F6E97",
x"8FC66F20",
x"90146F8C",
x"8FFC6FCD",
x"8F766FD4",
x"8E8A6FA0",
x"8D466F33",
x"8BC56E99",
x"8A256DE1",
x"88866D21",
x"87046C6C",
x"85B46BCF",
x"849A6B54",
x"83AE6AF3",
x"82D86A9A",
x"81F26A2E",
x"80CB698D",
x"7F386893",
x"7D0E6723",
x"7A346528",
x"769D62A4",
x"725B5FA7",
x"6D8F5C55",
x"687358DF",
x"634E5587",
x"5E6E5288",
x"5A1A501F",
x"56964E75",
x"540F4DA7",
x"529F4DB7",
x"52454E93",
x"52F15018",
x"54785213",
x"56AA5450",
x"594D5698",
x"5C2A58BC",
x"5F105A98",
x"61D65C18",
x"64655D35",
x"66AB5DF7",
x"68A65E6D",
x"6A595EAC",
x"6BCC5ECB",
x"6D0C5EDF",
x"6E215EF7",
x"6F175F1D",
x"6FF05F55",
x"70B25F9D",
x"715F5FEE",
x"71F76042",
x"7279608E",
x"72E860CF",
x"734260FA",
x"738E6110",
x"73CC610D",
x"740360F3",
x"743460C6",
x"74636088",
x"74906043",
x"74BD5FFA",
x"74E65FB7",
x"750A5F80",
x"75275F5D",
x"75385F58",
x"753C5F70",
x"75315FAB",
x"75176006",
x"74EF607C",
x"74BF6103",
x"748C6191",
x"745E621B",
x"743B6293",
x"742D62F2",
x"7438632E",
x"7460634B",
x"74A86349",
x"750C6332",
x"758A6315",
x"761E62FE",
x"76C162FC",
x"7770631A",
x"7826635C",
x"78DF63C6",
x"79986452",
x"7A4F64F3",
x"7B03659D",
x"7BAD663E",
x"7C4B66C6",
x"7CD66728",
x"7D4B675E",
x"7DA56762",
x"7DE6673E",
x"7E1366FD",
x"7E3466AE",
x"7E566665",
x"7E8A6632",
x"7EE26628",
x"7F696650",
x"802766B0",
x"81186741",
x"822F67FC",
x"835868CC",
x"846F69A3",
x"85566A65",
x"85E96B02",
x"86116B69",
x"85BE6B92",
x"84EF6B7A",
x"83B46B28",
x"82286AA8",
x"80726A0C",
x"7EBB6966",
x"7D2A68CC",
x"7BDC684B",
x"7AE867EF",
x"7A4F67B8",
x"7A0C67A8",
x"7A0967B1",
x"7A2F67C8",
x"7A6367DF",
x"7A9167E6",
x"7AAA67D2",
x"7AA867A0",
x"7A90674C",
x"7A6C66DF",
x"7A4B6660",
x"7A3B65DF",
x"7A476568",
x"7A706504",
x"7AB864BF",
x"7B13649B",
x"7B73649B",
x"7BC864BA",
x"7C0464EF",
x"7C1D6534",
x"7C0D657F",
x"7BD665C9",
x"7B81660E",
x"7B1D664B",
x"7AB7667D",
x"7A5D66A4",
x"7A1B66C2",
x"79F266D2",
x"79DC66D1",
x"79C966B8",
x"79A5667F",
x"7952661A",
x"78B26580",
x"77AB64A8",
x"762A6391",
x"7425623B",
x"71A360AF",
x"6EB55EFD",
x"6B7F5D38",
x"682A5B78",
x"64E959D9",
x"61EE586D",
x"5F62574A",
x"5D6B567A",
x"5C1D5601",
x"5B7D55DA",
x"5B8655FA",
x"5C23564F",
x"5D3656C4",
x"5E9E5749",
x"603D57CC",
x"61F55843",
x"63AB58AE",
x"6551590E",
x"66DC596D",
x"684459D7",
x"698A5A57",
x"6AAD5AFA",
x"6BAE5BBF",
x"6C915CA5",
x"6D595DA2",
x"6E0A5EA4",
x"6EA85F98",
x"6F3B606A",
x"6FCA610A",
x"705E616F",
x"70FD6198",
x"71B0618E",
x"72776163",
x"73536131",
x"743E6110",
x"752F611A",
x"761A6160",
x"76F561EC",
x"77B162BB",
x"784B63C1",
x"78BE64E3",
x"790E6606",
x"7941670A",
x"796367D1",
x"79836845",
x"79AE685B",
x"79F06813",
x"7A536779",
x"7ADE66A5",
x"7B8C65B7",
x"7C5964CE",
x"7D41640E",
x"7E386395",
x"7F376376",
x"803763BC",
x"81316469",
x"82276572",
x"831466C2",
x"83FD6841",
x"84DD69D1",
x"85B26B55",
x"86776CB4",
x"87226DD5",
x"87AB6EAB",
x"88036F30",
x"88246F61",
x"88076F47",
x"87B16EEB",
x"87276E5F",
x"867C6DB5",
x"85C46CFD",
x"85186C48",
x"84906BA3",
x"843F6B17",
x"84326AB0",
x"846C6A6D",
x"84E66A51",
x"85916A5B",
x"86566A86",
x"871D6ACE",
x"87C96B2B",
x"88496B96",
x"888D6C03",
x"88906C6B",
x"88586CC4",
x"87F06D06",
x"876D6D2B",
x"86E56D2E",
x"866C6D12",
x"86166CD4",
x"85ED6C7D",
x"85FA6C16",
x"863C6BA4",
x"86AA6B34",
x"87386ACB",
x"87D56A6F",
x"88706A21",
x"88F769E3",
x"895C69B1",
x"89916984",
x"89916959",
x"895D692D",
x"88F968FC",
x"887368CC",
x"87E268A3",
x"875F688A",
x"8707688E",
x"86F668BC",
x"87466920",
x"880869BE",
x"893F6A97",
x"8AE26BA7",
x"8CDA6CE2",
x"8F076E37",
x"91396F90",
x"934570DA",
x"94FE71FE",
x"964372E8",
x"96FD738D",
x"972573E5",
x"96C373EA",
x"95E9739D",
x"94AE7305",
x"932C7226",
x"917A7108",
x"8F9F6FB0",
x"8DA06E26",
x"8B706C70",
x"89036A96",
x"864668A0",
x"832F669A",
x"7FBC6493",
x"7BF7629B",
x"77FF60C2",
x"73F45F1A",
x"700D5DAF",
x"6C765C8B",
x"69625BB5",
x"66F25B29",
x"653D5AE1",
x"64475AD3",
x"64055AF3",
x"64615B32",
x"65385B84",
x"66655BE1",
x"67C55C42",
x"693A5CA5",
x"6AAD5D0B",
x"6C115D76",
x"6D605DEA",
x"6E9E5E6C",
x"6FCE5EFC",
x"70F65F9A",
x"72186042",
x"733B60F3",
x"745961A5",
x"75706255",
x"767C62FC",
x"77776398",
x"78606425",
x"793764A7",
x"79FF651B",
x"7ABE6586",
x"7B7C65E9",
x"7C3B6646",
x"7D0066A1",
x"7DC966F6",
x"7E906746",
x"7F466790",
x"7FDB67CE",
x"803E67FC",
x"805C6819",
x"80286820",
x"7F9B680E",
x"7EBA67E3",
x"7D8D679E",
x"7C2A6741",
x"7AAD66CE",
x"79346648",
x"77DD65B8",
x"76C46523",
x"75F96491",
x"7586640E",
x"756A63A3",
x"75A06358",
x"76116337",
x"76AE6342",
x"7760637D",
x"781463E3",
x"78BC6470",
x"794B6518",
x"79BE65CE",
x"7A136683",
x"7A4E6728",
x"7A7367B4",
x"7A8A681D",
x"7A976862",
x"7AA06886",
x"7AAB688D",
x"7ABD6880",
x"7AD9686C",
x"7B066859",
x"7B456851",
x"7B986856",
x"7BFF686D",
x"7C746894",
x"7CF268C5",
x"7D6A68FA",
x"7DD26931",
x"7E17695F",
x"7E306983",
x"7E0E699C",
x"7DB269A4",
x"7D2169A0",
x"7C696991",
x"7BA1697C",
x"7AE86961",
x"7A5D6945",
x"7A1E692D",
x"7A47691B",
x"7AE26914",
x"7BF26919",
x"7D69692A",
x"7F2B6947",
x"8111696B",
x"82F06993",
x"849B69B5",
x"85EC69CC",
x"86C669D1",
x"872169BF",
x"86FD6994",
x"86716952",
x"85A16903",
x"84B268B0",
x"83CF6865",
x"831F6831",
x"82BC681E",
x"82B56834",
x"83076873",
x"83A268D6",
x"846C6954",
x"854169DB",
x"85FD6A58",
x"86806ABA",
x"86B26AF3",
x"868A6AFA",
x"86076ACB",
x"853A6A6B",
x"843869E2",
x"8321693F",
x"82106894",
x"811D67ED",
x"80586758",
x"7FC166D8",
x"7F4F6670",
x"7EE96618",
x"7E7065C5",
x"7DC1656A",
x"7CB864F9",
x"7B3C6462",
x"7942639B",
x"76CB62A2",
x"73EA6177",
x"70C46022",
x"6D845EB2",
x"6A615D39",
x"678D5BCB",
x"653A5A7E",
x"63855969",
x"62835898",
x"62385819",
x"629757F3",
x"6386581F",
x"64E95898",
x"669B5952",
x"687D5A3B",
x"6A765B40",
x"6C725C53",
x"6E685D64",
x"70545E6C",
x"72355F67",
x"74106058",
x"75E66141",
x"77B7622D",
x"797D631E",
x"7B32641B",
x"7CCC6523",
x"7E41662E",
x"7F8C6732",
x"80AA6823",
x"819E68F0",
x"826F6991",
x"83286A00",
x"83D96A3A",
x"848A6A48",
x"85486A3A",
x"86146A20",
x"86F06A11",
x"87D06A1E",
x"88AE6A56",
x"897A6AC1",
x"8A2B6B5B",
x"8AB96C1C",
x"8B226CF3",
x"8B6C6DCF",
x"8BA16E9E",
x"8BD26F4F",
x"8C116FD9",
x"8C71703A",
x"8D037072",
x"8DCF708A",
x"8ED9708F",
x"9021708C",
x"919B708D",
x"933C709C",
x"94F670BB",
x"96B870EE",
x"98747130",
x"9A1C717C",
x"9BA571CE",
x"9D04721D",
x"9E2F7264",
x"9F1E729C",
x"9FC872C0",
x"A02472D0",
x"A02C72C8",
x"9FDF72AB",
x"9F3C727C",
x"9E49723E",
x"9D1471FB",
x"9BAF71BA",
x"9A317186",
x"98B67166",
x"97597165",
x"96337183",
x"955A71C3",
x"94DC721D",
x"94BF7288",
x"950072F8",
x"9592735E",
x"966373AC",
x"975973D5",
x"985873D4",
x"994573A6",
x"9A04734E",
x"9A8372D2",
x"9AB57243",
x"9A9471A7",
x"9A267110",
x"99767085",
x"9895700F",
x"97986FAE",
x"96956F65",
x"959B6F2E",
x"94B86EFF",
x"93EF6ED2",
x"93396E9C",
x"928D6E54",
x"91D86DF3",
x"91076D75",
x"900E6CD9",
x"8EE06C24",
x"8D7E6B5E",
x"8BF66A93",
x"8A5A69D4",
x"88CC6931",
x"876A68BB",
x"86586883",
x"85AB6890",
x"857468E2",
x"85B46975",
x"86566A37",
x"87416B14",
x"88496BF2",
x"89496CB3",
x"8A156D41",
x"8A906D8C",
x"8AA76D88",
x"8A586D3B",
x"89B16CB0",
x"88C96BF9",
x"87BE6B32",
x"86AC6A6F",
x"85AA69C1",
x"84C16932",
x"83EA68BF",
x"8314685B",
x"821D67EF",
x"80DD6762",
x"7F31669A",
x"7CFA6584",
x"7A2D6418",
x"76CE6258",
x"72F96058",
x"6EDF5E35",
x"6ABA5C17",
x"66D25A25",
x"63695887",
x"60BB5757",
x"5EEF56A8",
x"5E195678",
x"5E3356BA",
x"5F235757",
x"60BE582C",
x"62CE5917",
x"651759F8",
x"67695ABD",
x"69975B59",
x"6B895BCB",
x"6D315C1C",
x"6E945C60",
x"6FBF5CA8",
x"70C85D08",
x"71C25D8D",
x"72BE5E3D",
x"73C55F15",
x"74D9600D",
x"75F06113",
x"76FC6211",
x"77ED62F9",
x"78B263B7",
x"793C6441",
x"79866494",
x"798D64AF",
x"7958649D",
x"78F56466",
x"78706418",
x"77DC63C1",
x"7749636D",
x"76C56324",
x"765B62EF",
x"760F62CF",
x"75E862C6",
x"75E862D6",
x"761062FA",
x"7662632F",
x"76DC6374",
x"777D63C4",
x"7841641B",
x"79206477",
x"7A1164D6",
x"7B096532",
x"7BFA658D",
x"7CD865E2",
x"7D94662E",
x"7E2A6673",
x"7E9666B1",
x"7EDC66E9",
x"7F09671D",
x"7F2A6752",
x"7F51678A",
x"7F9367CB",
x"7FFF6817",
x"809E6873",
x"817968DF",
x"828A695C",
x"83C969E9",
x"85256A84",
x"868E6B27",
x"87EF6BCF",
x"89376C78",
x"8A586D1C",
x"8B4C6DB7",
x"8C106E47",
x"8CA56EC8",
x"8D146F3B",
x"8D636F9D",
x"8D9C6FEC",
x"8DC8702A",
x"8DE97054",
x"8E03706B",
x"8E12706E",
x"8E15705B",
x"8E047033",
x"8DD76FF6",
x"8D886FA4",
x"8D116F3E",
x"8C6A6EC4",
x"8B936E38",
x"8A8D6D9D",
x"895C6CF6",
x"880A6C45",
x"86A26B90",
x"85326ADE",
x"83C96A32",
x"82776997",
x"81466911",
x"804168A6",
x"7F706856",
x"7ED56828",
x"7E736819",
x"7E466826",
x"7E4F6849",
x"7E8B6880",
x"7EF968C4",
x"7F966913",
x"80636968",
x"815D69C5",
x"82806A2A",
x"83C46A96",
x"85186B09",
x"866F6B82",
x"87AF6BFA",
x"88C56C6B",
x"899B6CCD",
x"8A1F6D13",
x"8A496D38",
x"8A1B6D37",
x"899A6D0A",
x"88D96CB8",
x"87EC6C44",
x"86E76BB8",
x"85DF6B1D",
x"84D96A7C",
x"83DA69D6",
x"82D86930",
x"81BF6881",
x"807C67C1",
x"7EF666E5",
x"7D2065E5",
x"7AF364BB",
x"787A636C",
x"75CC6200",
x"7311608E",
x"70795F2E",
x"6E3B5E01",
x"6C8C5D28",
x"6B985CBD",
x"6B825CD6",
x"6C595D7B",
x"6E1E5EAC",
x"70BF605A",
x"741E6272",
x"781464D0",
x"7C77675B",
x"811A69ED",
x"85D56C70",
x"8A846ECE",
x"8F0E70F9",
x"935D72EF",
x"976474B3",
x"9B1B7648",
x"9E7B77BD",
x"A1847918",
x"A4367A64",
x"A6957BA5",
x"A8A67CDE",
x"AA717E0E",
x"ABFD7F2D",
x"AD53803A",
x"AE828129",
x"AF9681F1",
x"B09F828F",
x"B1A982FE",
x"B2C38342",
x"B3F78361",
x"B5518368",
x"B6D98368",
x"B88C8371",
x"BA6A8395",
x"BC6583E1",
x"BE6D8461",
x"C06A8512",
x"C24085EE",
x"C3D486E4",
x"C50C87DF",
x"C5D688C5",
x"C626897D",
x"C60489F7",
x"C57C8A28",
x"C4AC8A11",
x"C3B789C0",
x"C2C7894C",
x"C20488D3",
x"C18E8873",
x"C17B884A",
x"C1D6886D",
x"C29688E3",
x"C3A989A7",
x"C4F18AA8",
x"C6498BCB",
x"C7898CEA",
x"C8918DE3",
x"C93E8E96",
x"C97E8EE6",
x"C9428EC3",
x"C8878E2B",
x"C7518D22",
x"C5AC8BBC",
x"C3AA8A0E",
x"C1618836",
x"BEEB8652",
x"BC688481",
x"B9FA82DD",
x"B7C58181",
x"B5EA807E",
x"B4897FE0",
x"B3B97FB0",
x"B3877FEB",
x"B3F08088",
x"B4E18178",
x"B63C82A5",
x"B7D483F1",
x"B9778540",
x"BAEE8674",
x"BC0E8771",
x"BCAD8821",
x"BCBA8874",
x"BC2F8867",
x"BB1B87F9",
x"B9958733",
x"B7C38627",
x"B5C984E3",
x"B3C68378",
x"B1D481FB",
x"AFFB8077",
x"AE3D7EFC",
x"AC8E7D8F",
x"AAD77C3C",
x"A90A7B05",
x"A71279F2",
x"A4EE7903",
x"A2A1783C",
x"A03B779B",
x"9DDC771D",
x"9BA576C3",
x"99BB7681",
x"983E7652",
x"9745762F",
x"96D5760D",
x"96E675EA",
x"975D75BA",
x"9815757F",
x"98DC7533",
x"998174D5",
x"99D67467",
x"99B573E5",
x"990A7350",
x"97CF72A6",
x"960D71E6",
x"93DF7110",
x"91637026",
x"8EBF6F27",
x"8C146E14",
x"897A6CF3",
x"86FE6BC2",
x"84A16A82",
x"82526932",
x"7FFD67D1",
x"7D876656",
x"7AD564C2",
x"77D66310",
x"74806141",
x"70D95F59",
x"6CF95D62",
x"68FD5B67",
x"6510597E",
x"616257B8",
x"5E1C5626",
x"5B6554DD",
x"595A53E7",
x"58065349",
x"576C5304",
x"5782530F",
x"582E5363",
x"595A53ED",
x"5ADF549F",
x"5CA3556A",
x"5E835640",
x"60655715",
x"623357E3",
x"63DB58A4",
x"654F5955",
x"668A59F6",
x"67875A85",
x"684B5B05",
x"68D85B76",
x"69385BD5",
x"697B5C24",
x"69A85C61",
x"69D15C91",
x"6A005CB2",
x"6A3D5CCB",
x"6A8C5CDC",
x"6AEC5CEE",
x"6B5B5D06",
x"6BD15D28",
x"6C425D57",
x"6CAD5D95",
x"6D075DE0",
x"6D525E35",
x"6D915E8E",
x"6DC95EE4",
x"6E035F32",
x"6E455F70",
x"6E995F9D",
x"6EFD5FB7",
x"6F735FBE",
x"6FF35FB9",
x"70725FA9",
x"70E65F97",
x"71445F83",
x"71865F6E",
x"71AA5F59",
x"71B45F42",
x"71AD5F24",
x"71A15EFC",
x"71A05EC8",
x"71B75E8B",
x"71EC5E49",
x"72475E0B",
x"72C15DDD",
x"73535DC9",
x"73F05DD9",
x"74895E11",
x"750D5E76",
x"75755F00",
x"75BA5FA7",
x"75DB6059",
x"75DF610A",
x"75D261A5",
x"75BC6221",
x"75AE6272",
x"75AD6295",
x"75BC628E",
x"75DB6268",
x"76006229",
x"761E61E2",
x"762A619F",
x"7611616A",
x"75CC614B",
x"75566143",
x"74AF6158",
x"73E36184",
x"730261C5",
x"721D621A",
x"714C627E",
x"70A462EF",
x"70346368",
x"700763E5",
x"701D645F",
x"706D64CF",
x"70ED652A",
x"71876568",
x"7227657D",
x"72B86565",
x"7328651B",
x"736C64A3",
x"737C6403",
x"73596344",
x"730A6274",
x"729661A2",
x"720A60DC",
x"71726029",
x"70D85F92",
x"70455F17",
x"6FBF5EB5",
x"6F4C5E66",
x"6EEC5E24",
x"6EA35DE9",
x"6E6D5DB1",
x"6E4C5D77",
x"6E3F5D42",
x"6E425D10",
x"6E545CE7",
x"6E6D5CCB",
x"6E8A5CBC",
x"6EA45CBB",
x"6EB25CC2",
x"6EB05CCD",
x"6E995CD5",
x"6E695CD3",
x"6E215CC5",
x"6DC45CA4",
x"6D4F5C71",
x"6CC95C2F",
x"6C315BE0",
x"6B865B87",
x"6AC55B26",
x"69EB5AC0",
x"68F55A55",
x"67DF59E1",
x"66AB5969",
x"656158EA",
x"64075866",
x"62AE57E3",
x"61665766",
x"604256F7",
x"5F5456A1",
x"5EA9566A",
x"5E4A565A",
x"5E375677",
x"5E6E56BD",
x"5EE5572B",
x"5F9257BA",
x"60645861",
x"614F5915",
x"624F59CF",
x"635B5A81",
x"64725B26",
x"65975BBC",
x"66CF5C3D",
x"681E5CAB",
x"69855D0A",
x"6B025D5C",
x"6C965DAC",
x"6E375E00",
x"6FE05E60",
x"718A5ED9",
x"732B5F6E",
x"74C2602B",
x"764C610E",
x"77C9621A",
x"793C6345",
x"7AAA648A",
x"7C1465D6",
x"7D7A671A",
x"7EDC6845",
x"80316944",
x"81726A0C",
x"82936A91",
x"83846AD4",
x"843E6AD8",
x"84B16AA6",
x"84D86A4C",
x"84AF69DC",
x"843B6965",
x"838068F3",
x"828D6893",
x"81706848",
x"803F6817",
x"7F0E67FC",
x"7DF367F2",
x"7CFF67F0",
x"7C4467F5",
x"7BCE67F7",
x"7BA367F7",
x"7BC567F3",
x"7C2F67ED",
x"7CD967E9",
x"7DB567EB",
x"7EB467F5",
x"7FC2680E",
x"80D16837",
x"81CE686F",
x"82AF68B5",
x"836C6906",
x"83FC695E",
x"846069B7",
x"84976A0A",
x"84A76A56",
x"84946A96",
x"84696AC9",
x"842C6AF3",
x"83E96B14",
x"83A86B32",
x"83726B4F",
x"834E6B70",
x"83426B96",
x"83506BBF",
x"837C6BEC",
x"83BF6C19",
x"841A6C3E",
x"84866C5C",
x"84FB6C72",
x"85746C7F",
x"85ED6C89",
x"865F6C96",
x"86CB6CB0",
x"872F6CDF",
x"878E6D2A",
x"87EA6D93",
x"88436E19",
x"889B6EB4",
x"88EF6F57",
x"893B6FF0",
x"89797072",
x"89A270C7",
x"89B270E5",
x"89A270C3",
x"89727062",
x"89226FC8",
x"88BC6F02",
x"88496E23",
x"87D66D3E",
x"87746C6B",
x"87326BBA",
x"871D6B3A",
x"873F6AF7",
x"879D6AF5",
x"88346B31",
x"88FC6BA6",
x"89E76C4A",
x"8AE26D0C",
x"8BD86DDF",
x"8CB26EB1",
x"8D626F73",
x"8DD67017",
x"8E087094",
x"8DF970E2",
x"8DAC70FF",
x"8D3170EB",
x"8C9070AB",
x"8BD67044",
x"8B0A6FBA",
x"8A2B6F0F",
x"892B6E43",
x"87F66D52",
x"866F6C34",
x"84736ADC",
x"81E26941",
x"7EA46759",
x"7AAE6523",
x"7609629F",
x"70CE5FE0",
x"6B315CFB",
x"65755A0E",
x"5FE6573D",
x"5AD554AF",
x"568D5285",
x"534850D8",
x"512D4FBA",
x"50474F2D",
x"50864F29",
x"51C84F99",
x"53D55062",
x"566E5166",
x"594E5285",
x"5C3B53A6",
x"5F0454B6",
x"618C55AB",
x"63BD5681",
x"6597573F",
x"672357EE",
x"6870589A",
x"6990594F",
x"6A945A15",
x"6B895AF1",
x"6C765BE6",
x"6D5E5CEE",
x"6E415E04",
x"6F1D5F1E",
x"6FED6032",
x"70B16134",
x"7163621B",
x"720662DD",
x"72966374",
x"731863DD",
x"738C641A",
x"73F3642D",
x"744F641B",
x"74A363F2",
x"74F063BB",
x"753C6387",
x"75876362",
x"75D66353",
x"762A6365",
x"76836393",
x"76DC63DA",
x"7734642F",
x"77816486",
x"77BE64CC",
x"77E564F6",
x"77F264F7",
x"77E664CF",
x"77CB647F",
x"77AA6413",
x"7796639B",
x"779E632E",
x"77D862E0",
x"785162C8",
x"790D62F0",
x"7A106360",
x"7B4E6415",
x"7CB56504",
x"7E306617",
x"7FA0673A",
x"80EA684F",
x"81FC6942",
x"82C26A00",
x"83386A7F",
x"835D6ABD",
x"83416AC2",
x"82F36A9C",
x"828A6A5B",
x"821E6A16",
x"81C369DE",
x"818D69C4",
x"818369CE",
x"81AD6A03",
x"82076A5E",
x"82906AD7",
x"833B6B65",
x"83FF6BF9",
x"84D26C8C",
x"85AC6D10",
x"86846D83",
x"87566DE1",
x"881B6E26",
x"88D06E58",
x"89746E76",
x"8A016E85",
x"8A736E85",
x"8AC66E76",
x"8AF46E58",
x"8AF76E29",
x"8ACB6DE5",
x"8A696D8F",
x"89D06D21",
x"89016CA0",
x"88046C0D",
x"86E26B6B",
x"85A86AC2",
x"84696A19",
x"833C6979",
x"823568E9",
x"816A6875",
x"80EF6821",
x"80CC67F5",
x"810A67F2",
x"81A16819",
x"82866863",
x"83A268CB",
x"84DD6947",
x"861B69CB",
x"87426A4E",
x"883B6AC7",
x"88F96B2E",
x"89736B82",
x"89AE6BC5",
x"89B26BFA",
x"898D6C28",
x"894B6C54",
x"88F46C7F",
x"88916CA7",
x"881B6CC8",
x"87886CD5",
x"86C36CC1",
x"85BB6C7C",
x"84566BF9",
x"828A6B2E",
x"80516A19",
x"7DAF68BF",
x"7ABB6731",
x"77986583",
x"746F63D0",
x"71736239",
x"6ED460D8",
x"6CBB5FC2",
x"6B495F08",
x"6A935EB1",
x"6A975EB8",
x"6B495F12",
x"6C905FB2",
x"6E4B6084",
x"70526179",
x"72836280",
x"74C16390",
x"76F564A3",
x"791665B7",
x"7B2366CB",
x"7D1E67E0",
x"7F1468F6",
x"810C6A0A",
x"830D6B16",
x"851A6C13",
x"872E6CFA",
x"89416DC7",
x"8B466E72",
x"8D356F00",
x"8EFE6F73",
x"909E6FD5",
x"92117031",
x"93597093",
x"947D7103",
x"95847188",
x"96737221",
x"974F72CE",
x"98187382",
x"98CF7434",
x"996F74D5",
x"99F4755C",
x"9A6375C3",
x"9ABE7606",
x"9B0D7627",
x"9B5D7631",
x"9BC0762D",
x"9C437629",
x"9CF17630",
x"9DCF764E",
x"9EDC7686",
x"A00D76DE",
x"A14F7751",
x"A29177DA",
x"A3BB7871",
x"A4BB790F",
x"A58879AA",
x"A6217A3D",
x"A68A7AC0",
x"A6D37B32",
x"A7117B8F",
x"A7547BD9",
x"A7B57C0C",
x"A8397C2C",
x"A8E77C37",
x"A9B97C30",
x"AAA17C18",
x"AB8A7BF1",
x"AC5E7BC3",
x"AD087B93",
x"AD757B6A",
x"AD9C7B50",
x"AD7D7B50",
x"AD1B7B6D",
x"AC8A7BAD",
x"ABDC7C12",
x"AB2C7C96",
x"AA927D35",
x"AA247DE1",
x"A9EE7E8F",
x"A9FA7F33",
x"AA457FC3",
x"AAC38033",
x"AB648081",
x"AC1280A6",
x"ACB680A9",
x"AD3C808B",
x"AD958057",
x"ADB98014",
x"ADA67FCA",
x"AD647F85",
x"ACFE7F47",
x"AC807F18",
x"ABF67EF5",
x"AB687EDE",
x"AADA7ECF",
x"AA437EBD",
x"A9957EA3",
x"A8C07E78",
x"A7B07E2F",
x"A6567DC3",
x"A4A57D2C",
x"A29F7C6A",
x"A04F7B7C",
x"9DCF7A6D",
x"9B3C7946",
x"98C07819",
x"968476F8",
x"94AA75F5",
x"934C751F",
x"927A7483",
x"92347425",
x"92697400",
x"9300740D",
x"93D5743E",
x"94BF7480",
x"959F74C4",
x"965674FB",
x"96D3751F",
x"9712752F",
x"971E752F",
x"9706752C",
x"96E2752F",
x"96C97543",
x"96CB756B",
x"96EC75A5",
x"972275E2",
x"9758760C",
x"97627608",
x"971175B6",
x"963274F9",
x"949573C0",
x"921D71FF",
x"8EB96FBD",
x"8A746D0C",
x"85716A0D",
x"7FEA66E9",
x"7A2A63CC",
x"748360E4",
x"6F485E56",
x"6AC45C3D",
x"672B5AA9",
x"649E599F",
x"63235915",
x"62A858FB",
x"6309593C",
x"641359BF",
x"65905A6D",
x"674B5B35",
x"69195C06",
x"6AD75CD5",
x"6C725D9C",
x"6DE25E5A",
x"6F2D5F0E",
x"70595FB9",
x"7175605D",
x"728760FC",
x"739B6194",
x"74B46228",
x"75D162B8",
x"76EF6342",
x"780A63C4",
x"791D643F",
x"7A2464B1",
x"7B1B6517",
x"7BFF656F",
x"7CCE65BA",
x"7D8365F3",
x"7E1A661A",
x"7E8B6630",
x"7ED36634",
x"7EEC6627",
x"7ED36609",
x"7E8965DE",
x"7E1665A5",
x"7D836563",
x"7CE0651A",
x"7C3E64CE",
x"7BAE6483",
x"7B3C643C",
x"7AF46401",
x"7AD663D3",
x"7ADF63B5",
x"7B0363AA",
x"7B3463AF",
x"7B6063C5",
x"7B7A63E8",
x"7B776415",
x"7B566448",
x"7B186481",
x"7ACB64BC",
x"7A7C64FF",
x"7A416549",
x"7A2865A0",
x"7A416604",
x"7A906679",
x"7B1466FD",
x"7BBF678A",
x"7C83681A",
x"7D48689E",
x"7DF7690D",
x"7E80695B",
x"7ED2697F",
x"7EE76975",
x"7EC5693E",
x"7E7368E5",
x"7DFF6875",
x"7D7A6800",
x"7CF66799",
x"7C80674C",
x"7C216727",
x"7BDB672B",
x"7BAA6758",
x"7B89679E",
x"7B6D67F0",
x"7B4F6838",
x"7B276863",
x"7AEF6862",
x"7AA76827",
x"7A5367B2",
x"79F96709",
x"799E6637",
x"7949654F",
x"79006466",
x"78BF6390",
x"788762DC",
x"78536255",
x"781A61FE",
x"77D361D5",
x"777961CF",
x"770761DF",
x"767C61F6",
x"75D96209",
x"7527620D",
x"746D61FC",
x"73B761D8",
x"730E61A5",
x"727A616A",
x"7202612F",
x"71A360FE",
x"715B60D9",
x"712460C1",
x"70F360B4",
x"70BE60A9",
x"707C609A",
x"7027607D",
x"6FB8604C",
x"6F326003",
x"6E965F9F",
x"6DE95F25",
x"6D345E9A",
x"6C7A5E03",
x"6BC25D69",
x"6B0E5CD3",
x"6A5E5C43",
x"69B05BBD",
x"68FD5B3F",
x"68445AC5",
x"677C5A4A",
x"66A459CA",
x"65B75942",
x"64B858AE",
x"63A8580B",
x"6290575C",
x"617256A1",
x"605A55E0",
x"5F4B551E",
x"5E525460",
x"5D7353AD",
x"5CB6530C",
x"5C205285",
x"5BB4521F",
x"5B7951DD",
x"5B7251C7",
x"5BA051DE",
x"5C065225",
x"5CA0529B",
x"5D6F533C",
x"5E6B5405",
x"5F8C54EE",
x"60CB55F3",
x"621D5707",
x"63795824",
x"64D45942",
x"66265A59",
x"67695B61",
x"689A5C56",
x"69B55D31",
x"6ABB5DED",
x"6BAA5E8A",
x"6C845F07",
x"6D485F64",
x"6DF65FA7",
x"6E8D5FD6",
x"6F0D5FF9",
x"6F766018",
x"6FC8603E",
x"70056070",
x"703160B4",
x"7051610A",
x"706C6173",
x"708961EC",
x"70B0626D",
x"70E862F3",
x"71356373",
x"719D63EA",
x"72216453",
x"72C264AB",
x"737C64ED",
x"7448651A",
x"75216531",
x"75FD652F",
x"76D16517",
x"779164E5",
x"7838649E",
x"78BC6446",
x"791D63E5",
x"795B6383",
x"797D6331",
x"799062FC",
x"79A262F3",
x"79C76324",
x"7A0C6395",
x"7A80644B",
x"7B2F6541",
x"7C1D666C",
x"7D4467BA",
x"7E976917",
x"800A6A6D",
x"81846BA7",
x"82F36CB5",
x"84446D8C",
x"85676E26",
x"86556E85",
x"870B6EB3",
x"87916EB8",
x"87F36EA4",
x"883E6E83",
x"88836E61",
x"88D06E44",
x"89356E34",
x"89B56E31",
x"8A536E38",
x"8B0B6E4A",
x"8BD86E61",
x"8CAB6E79",
x"8D7B6E94",
x"8E3B6EB0",
x"8EDF6ECE",
x"8F5F6EF0",
x"8FB76F19",
x"8FE26F45",
x"8FE26F76",
x"8FB86FA7",
x"8F676FD2",
x"8EF36FF0",
x"8E5C6FF8",
x"8DA46FDF",
x"8CCC6FA0",
x"8BD56F34",
x"8AC16E99",
x"89936DCF",
x"88506CE1",
x"87036BD7",
x"85B66ABD",
x"847C69A6",
x"836068A1",
x"827467BE",
x"81C26709",
x"8151668B",
x"81206645",
x"81276635",
x"81586650",
x"819B668A",
x"81D966D1",
x"81FA6713",
x"81E86741",
x"81946749",
x"80F96725",
x"801D66CF",
x"7F0B664C",
x"7DDB65A5",
x"7CA364E6",
x"7B7A6423",
x"7A73636D",
x"799862D6",
x"78EC626D",
x"78626237",
x"77E66234",
x"7762625D",
x"76BE62A4",
x"75E062F4",
x"74C16338",
x"735B6356",
x"71BA633C",
x"6FF362DF",
x"6E256239",
x"6C756150",
x"6B066035",
x"69F35F00",
x"69565DCB",
x"69355CB8",
x"69905BE1",
x"6A565B61",
x"6B725B45",
x"6CC75B92",
x"6E3A5C45",
x"6FAE5D49",
x"71105E8B",
x"72525FEC",
x"736F614E",
x"74686297",
x"754263AF",
x"7609648B",
x"76C66525",
x"77876583",
x"785265B1",
x"793165C2",
x"7A2865CF",
x"7B3965EC",
x"7C656628",
x"7DA76690",
x"7EFF6725",
x"806367E2",
x"81CF68B7",
x"83376993",
x"84916A5F",
x"85D36B0A",
x"86F66B86",
x"87F06BCE",
x"88BE6BE2",
x"895D6BCE",
x"89D36BA4",
x"8A216B76",
x"8A4E6B57",
x"8A606B57",
x"8A5F6B7C",
x"8A4C6BC7",
x"8A2C6C31",
x"8A046CAB",
x"89D36D27",
x"899F6D93",
x"896F6DE6",
x"89486E17",
x"89376E2A",
x"89456E24",
x"897E6E10",
x"89E96DFC",
x"8A896DF0",
x"8B5F6DF6",
x"8C626E0F",
x"8D886E3B",
x"8EC56E73",
x"90066EB3",
x"913C6EF5",
x"925D6F35",
x"935F6F78",
x"943B6FC1",
x"94ED7017",
x"95777083",
x"95D97106",
x"961271A1",
x"9624724D",
x"961072F6",
x"95D3738F",
x"95737400",
x"94F17434",
x"9457741F",
x"93AE73B6",
x"930472FC",
x"926471FE",
x"91DD70CD",
x"91776F82",
x"91346E37",
x"91136D03",
x"910B6BF9",
x"91106B24",
x"91106A86",
x"90F96A1A",
x"90BB69D5",
x"904869AB",
x"8F9D698E",
x"8EB56973",
x"8D9B694F",
x"8C566923",
x"8AF968EF",
x"899068BA",
x"882B688A",
x"86D9686C",
x"85A26862",
x"848A6870",
x"83936896",
x"82BB68CB",
x"82006906",
x"815B693E",
x"80C96965",
x"804B6973",
x"7FDC695F",
x"7F7F692B",
x"7F3468D8",
x"7EFC686C",
x"7ED567F3",
x"7EBF6776",
x"7EB266FD",
x"7EAA6690",
x"7E9D662D",
x"7E8165D5",
x"7E526581",
x"7E06652D",
x"7D9D64D0",
x"7D176468",
x"7C7963F4",
x"7BC8637A",
x"7B0D6303",
x"7A4E6298",
x"79906243",
x"78D5620A",
x"781761ED",
x"775161E3",
x"767261E0",
x"756A61CE",
x"742A6193",
x"729E611B",
x"70B86050",
x"6E705F29",
x"6BC55DA8",
x"68C25BD7",
x"657959CF",
x"620657AF",
x"5E8F559E",
x"5B3D53BF",
x"583D5236",
x"55B85118",
x"53D45072",
x"52AB5044",
x"524B5084",
x"52B4511B",
x"53D851EE",
x"559C52E1",
x"57DB53D7",
x"5A6954BA",
x"5D1A557B",
x"5FC25611",
x"623B567B",
x"646956BF",
x"663A56E9",
x"67A55702",
x"68B05719",
x"695F573A",
x"69C5576B",
x"69F357B2",
x"69FD580F",
x"69F25881",
x"69DF5901",
x"69CF598A",
x"69C85A14",
x"69CB5A95",
x"69D85B07",
x"69EB5B60",
x"6A035B9A",
x"6A1D5BB2",
x"6A385BA5",
x"6A545B77",
x"6A765B2B",
x"6AA05ACC",
x"6AD95A64",
x"6B235A04",
x"6B8059B8",
x"6BEF598E",
x"6C6C598F",
x"6CEC59C3",
x"6D635A28",
x"6DC55AB9",
x"6E045B6B",
x"6E165C31",
x"6DF55CF7",
x"6D9E5DAF",
x"6D1D5E48",
x"6C7A5EB9",
x"6BCB5EFE",
x"6B265F17",
x"6A9E5F08",
x"6A4E5EE3",
x"6A415EB1",
x"6A835E83",
x"6B165E64",
x"6BF25E62",
x"6D075E7E",
x"6E445EBB",
x"6F8D5F10",
x"70C85F74",
x"71DD5FDC",
x"72B5603C",
x"73416088",
x"737360B9",
x"734C60CC",
x"72CF60BF",
x"7207609A",
x"71096062",
x"6FE6601F",
x"6EBA5FDC",
x"6D9D5F9E",
x"6CA65F6E",
x"6BE85F4D",
x"6B725F3E",
x"6B495F3F",
x"6B725F4F",
x"6BE15F6A",
x"6C8A5F91",
x"6D5C5FBF",
x"6E425FF3",
x"6F28602B",
x"6FFC6063",
x"70AE6097",
x"713460C3",
x"718A60E6",
x"71B260F9",
x"71B160FA",
x"718D60E7",
x"715260C2",
x"7109608D",
x"70B46048",
x"70595FF7",
x"6FF95F9D",
x"6F8F5F3B",
x"6F195ED0",
x"6E915E5A",
x"6DF85DDA",
x"6D4B5D4C",
x"6C8D5CB1",
x"6BC85C0A",
x"6B025B5D",
x"6A485AB5",
x"69A65A1A",
x"69245998",
x"68CA5939",
x"68995905",
x"68915900",
x"68AA5925",
x"68D95970",
x"691159D3",
x"69445A3F",
x"69625AA8",
x"69625AFD",
x"693C5B36",
x"68F05B4B",
x"687D5B3C",
x"67EB5B0B",
x"67445AC0",
x"66915A64",
x"65DC59FE",
x"65305998",
x"648C5936",
x"63F058DD",
x"6359588E",
x"62BB5847",
x"620C5807",
x"614057CC",
x"604E5795",
x"5F355761",
x"5DF65732",
x"5C9E5707",
x"5B4056E1",
x"59F356C2",
x"58D256A9",
x"57FB5697",
x"5782568A",
x"5779567E",
x"57E85677",
x"58C85674",
x"5A105677",
x"5BA65681",
x"5D6C569B",
x"5F4456C6",
x"61105708",
x"62B45763",
x"641E57D6",
x"6542585D",
x"661C58F5",
x"66AE5995",
x"67045A33",
x"672A5AC7",
x"672E5B4B",
x"67205BB6",
x"670A5C0B",
x"66F85C49",
x"66EE5C71",
x"66EF5C8A",
x"67005C95",
x"671E5C97",
x"67485C8E",
x"677F5C7E",
x"67C15C66",
x"680A5C43",
x"685E5C1B",
x"68BA5BF0",
x"691D5BC9",
x"69875BAF",
x"69F55BA9",
x"6A635BBF",
x"6ACC5BF4",
x"6B275C46",
x"6B6F5CB1",
x"6B985D25",
x"6BA15D94",
x"6B835DED",
x"6B3F5E22",
x"6ADE5E29",
x"6A685E01",
x"69EF5DAE",
x"69855D3D",
x"69385CC5",
x"691A5C57",
x"69325C08",
x"69805BE7",
x"69FF5BFB",
x"6A9D5C42",
x"6B475CB2",
x"6BE65D3B",
x"6C665DC8",
x"6CB45E45",
x"6CC85EA1",
x"6C9E5ED3",
x"6C415EDA",
x"6BBA5EB9",
x"6B1D5E7D",
x"6A7C5E31",
x"69E85DE4",
x"696D5DA4",
x"69145D74",
x"68DB5D59",
x"68BE5D4F",
x"68B85D52",
x"68C05D5A",
x"68CE5D62",
x"68DF5D67",
x"68EF5D6A",
x"69025D6E",
x"691A5D7A",
x"693C5D92",
x"696D5DBC",
x"69AE5DFA",
x"6A025E48",
x"6A635E9F",
x"6AD25EF7",
x"6B475F43",
x"6BBB5F7D",
x"6C2B5F9B",
x"6C935F9D",
x"6CEF5F86",
x"6D3E5F5C",
x"6D845F29",
x"6DC45EF8",
x"6DFD5ED2",
x"6E335EB9",
x"6E655EAF",
x"6E935EB1",
x"6EB75EB3",
x"6ECB5EAC",
x"6EC55E90",
x"6E9D5E56",
x"6E4B5DFA",
x"6DCB5D7D",
x"6D1B5CE4",
x"6C425C3D",
x"6B4B5B97",
x"6A425AFE",
x"69405A82",
x"68545A2E",
x"67965A07",
x"67145A0D",
x"66D95A3C",
x"66E85A8D",
x"67375AF4",
x"67BA5B64",
x"685E5BD5",
x"690A5C39",
x"69A75C8E",
x"6A1C5CCF",
x"6A585CF6",
x"6A4A5D02",
x"69EC5CF4",
x"693A5CCB",
x"68345C81",
x"66E45C1A",
x"654F5B92",
x"63855AEE",
x"61905A30",
x"5F83595F",
x"5D705882",
x"5B6E57A8",
x"599056D9",
x"57EE5621",
x"569C5588",
x"55AC5516",
x"552C54CD",
x"552054AB",
x"558C54AC",
x"566554CA",
x"57A05501",
x"5929554D",
x"5AEC55A9",
x"5CD15618",
x"5EC55699",
x"60B55730",
x"629457E0",
x"645758A8",
x"65F85985",
x"67755A71",
x"68CB5B63",
x"69FC5C4F",
x"6B095D29",
x"6BF25DE9",
x"6CB75E86",
x"6D5B5EFC",
x"6DDC5F4C",
x"6E3B5F7A",
x"6E795F8B",
x"6E975F88",
x"6E975F76",
x"6E7D5F5A",
x"6E4C5F38",
x"6E0A5F10",
x"6DBF5EE0",
x"6D735EAC",
x"6D315E71",
x"6D035E36",
x"6CF25DFD",
x"6D065DCF",
x"6D445DB3",
x"6DAB5DAF",
x"6E3B5DCB",
x"6EE95E01",
x"6FA85E53",
x"70695EB3",
x"711A5F1B",
x"71AD5F7C",
x"72145FC8",
x"72495FF7",
x"72486007",
x"72145FF6",
x"71BA5FCC",
x"71425F94",
x"70BF5F5A",
x"703E5F2E",
x"6FCB5F1A",
x"6F705F27",
x"6F325F56",
x"6F135FA9",
x"6F106018",
x"6F25609A",
x"6F516122",
x"6F8F61A9",
x"6FE06227",
x"704A6293",
x"70CB62EF",
x"716B6339",
x"722B6376",
x"731063AA",
x"741163D6",
x"75286400",
x"76486425",
x"775E6446",
x"78596460",
x"7927646F",
x"79BA6470",
x"7A096460",
x"7A11643F",
x"79D8640E",
x"796863CF",
x"78CE6387",
x"781D633C",
x"776562F3",
x"76B162B2",
x"760F627D",
x"75806259",
x"75096248",
x"74A86249",
x"745B625C",
x"741E627A",
x"73F062A1",
x"73D162C8",
x"73BE62E6",
x"73BA62F6",
x"73C162EF",
x"73D262CC",
x"73E6628B",
x"73F9622D",
x"740261B4",
x"73F96125",
x"73DB6088",
x"73A45FE9",
x"73595F50",
x"72FF5EC5",
x"72A05E50",
x"72455DF8",
x"71FA5DC1",
x"71C45DA9",
x"71A65DB2",
x"719C5DDA",
x"71A35E1C",
x"71AE5E77",
x"71B55EE2",
x"71B05F58",
x"71965FD0",
x"71626043",
x"711660A7",
x"70B160F0",
x"703A6117",
x"6FAD6110",
x"6F0C60D3",
x"6E52605D",
x"6D765FAC",
x"6C6F5EC2",
x"6B315DA2",
x"69B55C57",
x"67F95AF0",
x"6600597B",
x"63D7580A",
x"619156AF",
x"5F4D557D",
x"5D2A5482",
x"5B4B53CC",
x"59CF5363",
x"58D2534A",
x"5866537F",
x"589653FD",
x"595F54B8",
x"5AB755A2",
x"5C8C56AE",
x"5EC457C7",
x"614258E4",
x"63EB59F7",
x"66A15AF6",
x"694E5BDF",
x"6BDB5CB1",
x"6E3B5D6D",
x"70635E1A",
x"72525EBD",
x"74065F5D",
x"75835FFD",
x"76CF609F",
x"77F56143",
x"78F761E8",
x"79DF6286",
x"7AAF6317",
x"7B686395",
x"7C0763FC",
x"7C8A6445",
x"7CEA6470",
x"7D256480",
x"7D356477",
x"7D1A645D",
x"7CD96439",
x"7C7A6415",
x"7C0763F6",
x"7B8E63DF",
x"7B2063D2",
x"7AC563CE",
x"7A8963CE",
x"7A6F63CC",
x"7A7663C5",
x"7A9863B4",
x"7AC96398",
x"7AFE6376",
x"7B2D6350",
x"7B4B632F",
x"7B58631D",
x"7B53631F",
x"7B48633F",
x"7B3F637D",
x"7B4963DA",
x"7B706453",
x"7BBC64DE",
x"7C2E6570",
x"7CBE6600",
x"7D606683",
x"7E0066EF",
x"7E86673E",
x"7EDD676D",
x"7EF7677C",
x"7EC8676B",
x"7E52673F",
x"7DA06701",
x"7CC566B8",
x"7BDE6670",
x"7B036631",
x"7A526606",
x"79E265FA",
x"79BE6613",
x"79E96653",
x"7A5D66BC",
x"7B096746",
x"7BD667E6",
x"7CAE688A",
x"7D756921",
x"7E1A6996",
x"7E9169D6",
x"7ED369D8",
x"7EE36994",
x"7ECB690D",
x"7E97684E",
x"7E536769",
x"7E0D6675",
x"7DCB658A",
x"7D9164BE",
x"7D5E6423",
x"7D2D63BE",
x"7CF66391",
x"7CB26394",
x"7C5F63B9",
x"7BF663ED",
x"7B7A641D",
x"7AF06438",
x"7A5B6434",
x"79C4640B",
x"792E63BF",
x"789E6359",
x"781662E3",
x"7794626D",
x"77166203",
x"769961B1",
x"7619617D",
x"7597616C",
x"7517617E",
x"749E61B1",
x"743461FD",
x"73E3625D",
x"73B762CB",
x"73B4633E",
x"73DC63AD",
x"74316411",
x"74AB6463",
x"753C649B",
x"75DB64B5",
x"767264AB",
x"76F5647F",
x"7753642F",
x"778463C6",
x"77806349",
x"774262C4",
x"76C8623C",
x"761161BE",
x"7520614B",
x"73F060E2",
x"72876081",
x"70E3601F",
x"6F0A5FB2",
x"6D035F31",
x"6AD95E92",
x"689D5DD5",
x"66665CFA",
x"644B5C0B",
x"62655B14",
x"60CE5A28",
x"5F975955",
x"5ECE58A8",
x"5E78582F",
x"5E9057EB",
x"5F0C57DD",
x"5FDC57FD",
x"60EB5840",
x"6226589C",
x"63795907",
x"64D75978",
x"663759EA",
x"67915A5C",
x"68E35AD0",
x"6A2D5B4B",
x"6B6C5BCC",
x"6CA05C55",
x"6DC45CE4",
x"6ED55D74",
x"6FCC5E00",
x"70A85E80",
x"71685EF0",
x"720A5F4D",
x"72965F9D",
x"73115FE3",
x"7383602B",
x"73F4607D",
x"746C60E3",
x"74E96162",
x"756F61FA",
x"75F762A5",
x"76806358",
x"77006404",
x"7775649B",
x"77DD6510",
x"783C6558",
x"78966573",
x"78F26566",
x"7959653B",
x"79D16501",
x"7A5D64CC",
x"7AFE64A8",
x"7BB164A5",
x"7C6A64CB",
x"7D256518",
x"7DD6658E",
x"7E776624",
x"7F0766D1",
x"7F876789",
x"7FFD6845",
x"80736900",
x"80EF69B2",
x"81776A5B",
x"82136AF7",
x"82B96B86",
x"83666C03",
x"840B6C6F",
x"849B6CC5",
x"850A6D03",
x"854B6D28",
x"855B6D35",
x"853F6D2B",
x"85036D12",
x"84B46CEB",
x"84666CBE",
x"842E6C93",
x"841B6C6C",
x"84386C4B",
x"84846C31",
x"84F96C1C",
x"85896C04",
x"861E6BE6",
x"86A46BBD",
x"87036B84",
x"872B6B3D",
x"87106AE6",
x"86AF6A83",
x"86106A1C",
x"853C69B2",
x"8445694E",
x"833F68F5",
x"823E68A7",
x"814F6869",
x"8080683A",
x"7FD56819",
x"7F4B6801",
x"7EDD67F5",
x"7E8367ED",
x"7E2E67EB",
x"7DD367E9",
x"7D6D67E6",
x"7CF767E2",
x"7C7367D9",
x"7BE367CC",
x"7B5367B8",
x"7ACE679B",
x"7A5D6779",
x"7A0D674F",
x"79E06720",
x"79DB66F0",
x"79F766C4",
x"7A2E669B",
x"7A74667C",
x"7ABE6663",
x"7AFC6652",
x"7B256641",
x"7B31662E",
x"7B186611",
x"7ADF65E8",
x"7A8365AD",
x"7A0D6560",
x"79836507",
x"78EB64A7",
x"78496446",
x"77A063EA",
x"76EC6398",
x"762A634E",
x"754F6306",
x"745162B4",
x"73256249",
x"71C161B5",
x"701E60E9",
x"6E3E5FDA",
x"6C235E86",
x"69DC5CF4",
x"677F5B36",
x"65245966",
x"62EC57A2",
x"60F5560F",
x"5F5C54C9",
x"5E3D53E8",
x"5DA4537D",
x"5D9C5389",
x"5E245404",
x"5F3154DC",
x"60B355F8",
x"6293573D",
x"64BA5894",
x"671159E6",
x"69865B28",
x"6C075C52",
x"6E8A5D6A",
x"71075E74",
x"73795F7D",
x"75D9608E",
x"782261AD",
x"7A5162DA",
x"7C596418",
x"7E37655E",
x"7FE066A3",
x"815267DB",
x"828D6901",
x"83956A11",
x"84746B07",
x"85386BE8",
x"85EF6CB5",
x"86A46D78",
x"87656E34",
x"88376EEB",
x"89156F9C",
x"89FD7043",
x"8ADD70D7",
x"8BAA714E",
x"8C4F71A3",
x"8CC271CA",
x"8CF971C1",
x"8CF17186",
x"8CB1711D",
x"8C45708F",
x"8BBC6FE2",
x"8B2F6F24",
x"8AB46E63",
x"8A5D6DAE",
x"8A3F6D10",
x"8A626C96",
x"8ACC6C47",
x"8B7A6C2B",
x"8C626C45",
x"8D706C94",
x"8E926D12",
x"8FAF6DB0",
x"90B16E62",
x"91836F16",
x"92156FB7",
x"925F7034",
x"9260707F",
x"9222708F",
x"91B27064",
x"91257003",
x"90916F7F",
x"900A6EE8",
x"8FA26E57",
x"8F666DE3",
x"8F586DA3",
x"8F736D9E",
x"8FAE6DE1",
x"8FFA6E65",
x"90466F1E",
x"90836FFE",
x"90A470E8",
x"90A171C8",
x"907C7286",
x"9038730D",
x"8FDC7354",
x"8F727354",
x"8F077312",
x"8EA27299",
x"8E4B71FE",
x"8E067155",
x"8DD270B7",
x"8DAF7039",
x"8D9B6FE9",
x"8D956FD4",
x"8D9A6FF6",
x"8DA7704A",
x"8DBB70BE",
x"8DD67140",
x"8DF371B9",
x"8E127213",
x"8E2F7241",
x"8E46723D",
x"8E577209",
x"8E6271AF",
x"8E67713E",
x"8E6D70D1",
x"8E7A707C",
x"8E977052",
x"8ECF705F",
x"8F2570AA",
x"8F9D712E",
x"903571DC",
x"90E372A3",
x"919A736B",
x"9245741C",
x"92D2749F",
x"932E74E2",
x"934974DC",
x"931E7489",
x"92AC73EC",
x"92007312",
x"91287206",
x"903C70DC",
x"8F506FA9",
x"8E776E7C",
x"8DB96D65",
x"8D146C69",
x"8C796B8D",
x"8BCB6AC9",
x"8AE76A13",
x"89A26959",
x"87D56889",
x"855D678E",
x"822A6656",
x"7E3764D8",
x"799A630B",
x"747860F7",
x"6F0A5EA9",
x"69965C39",
x"646259C3",
x"5FB7576A",
x"5BD25550",
x"58E15393",
x"56FF524C",
x"562E5187",
x"5661514A",
x"5772518F",
x"59315246",
x"5B685358",
x"5DDE54A9",
x"6061561F",
x"62C5579C",
x"64F3590B",
x"66DC5A5D",
x"68805B8A",
x"69EC5C8E",
x"6B345D6E",
x"6C6F5E36",
x"6DB35EEE",
x"6F115FA2",
x"7094605C",
x"723E611F",
x"740661EA",
x"75DC62B9",
x"77AE6380",
x"79636432",
x"7AE864C5",
x"7C2B652D",
x"7D246562",
x"7DCC6566",
x"7E2B653E",
x"7E4B64F6",
x"7E3C64A0",
x"7E13644C",
x"7DDF6411",
x"7DB463FD",
x"7D9D641B",
x"7DA06470",
x"7DBE64FA",
x"7DF665B1",
x"7E416683",
x"7E946763",
x"7EE9683E",
x"7F376903",
x"7F7C69A7",
x"7FB76A24",
x"7FEF6A76",
x"802B6AA4",
x"80746AB1",
x"80D56AAA",
x"81566A99",
x"81FC6A87",
x"82C86A7F",
x"83B56A84",
x"84BC6A9C",
x"85CF6AC5",
x"86DF6B03",
x"87DF6B4E",
x"88BE6BA6",
x"89706C06",
x"89ED6C69",
x"8A2F6CCB",
x"8A386D2A",
x"8A0A6D7D",
x"89AB6DC5",
x"89226DFC",
x"887D6E1E",
x"87C36E2A",
x"87036E1D",
x"86426DF9",
x"858D6DBE",
x"84E96D72",
x"845D6D1A",
x"83EC6CBD",
x"83986C63",
x"835F6C16",
x"833C6BD5",
x"832D6BA7",
x"83276B8A",
x"83246B76",
x"831B6B66",
x"83096B4E",
x"82E66B23",
x"82AE6ADB",
x"825F6A6F",
x"81FA69DB",
x"81806921",
x"80F3684B",
x"80566763",
x"7FAB6677",
x"7EF96598",
x"7E3F64D5",
x"7D866438",
x"7CCE63C9",
x"7C1B638B",
x"7B76637A",
x"7AE26393",
x"7A6563CB",
x"7A02641D",
x"79C16480",
x"79A464EF",
x"79AF6568",
x"79E565E8",
x"7A42666C",
x"7AC866F5",
x"7B6F677D",
x"7C3267FF",
x"7D0A6872",
x"7DEC68CC",
x"7ECE6909",
x"7FA76920",
x"806D690E",
x"811B68D8",
x"81A56881",
x"82066816",
x"823767A0",
x"822D672B",
x"81DF66BF",
x"8142665E",
x"804B6603",
x"7EEB65A7",
x"7D19653A",
x"7ACF64AE",
x"780D63F2",
x"74DE62FE",
x"715361CE",
x"6D896064",
x"69A35ED0",
x"65CF5D24",
x"623A5B78",
x"5F0F59E6",
x"5C735885",
x"5A825767",
x"5948569B",
x"58C55621",
x"58EB55F5",
x"599D560F",
x"5ABD5661",
x"5C2156D7",
x"5DA75763",
x"5F3157F3",
x"60A4587A",
x"61F358F1",
x"63145950",
x"640A5998",
x"64D559C6",
x"657F59E0",
x"660C59EB",
x"668059F1",
x"66E459FD",
x"67335A15",
x"67755A47",
x"67A95A9B",
x"67D55B17",
x"68005BBC",
x"68345C87",
x"68785D6E",
x"68D25E64",
x"694B5F59",
x"69E2603B",
x"6A9460F7",
x"6B5B6180",
x"6C2761CF",
x"6CEC61E0",
x"6D9D61B9",
x"6E306164",
x"6E9A60F3",
x"6EDB6073",
x"6EF35FF7",
x"6EEB5F8E",
x"6EC85F45",
x"6E975F21",
x"6E635F22",
x"6E345F49",
x"6E135F8D",
x"6E035FE4",
x"6E0A6049",
x"6E2860B2",
x"6E606115",
x"6EB1616D",
x"6F1D61B4",
x"6FA161E8",
x"703C6206",
x"70EC620E",
x"71AA6204",
x"726D61EA",
x"732D61C3",
x"73DF619A",
x"74786173",
x"74F06158",
x"75426150",
x"756D6162",
x"75756190",
x"756061DA",
x"753F623E",
x"751E62B1",
x"750E632A",
x"75206398",
x"755F63F4",
x"75D16434",
x"76776452",
x"774C644F",
x"78426434",
x"7949640A",
x"7A4B63E5",
x"7B3163D2",
x"7BE963E2",
x"7C63641D",
x"7C976486",
x"7C846517",
x"7C3265C5",
x"7BAD667F",
x"7B09672D",
x"7A5967BA",
x"79B46817",
x"79286838",
x"78C46819",
x"788A67BE",
x"787A6734",
x"788D668A",
x"78B865D5",
x"78F06521",
x"792B6480",
x"796363F9",
x"7998638B",
x"79CC6337",
x"7A0762F3",
x"7A4F62BC",
x"7AAB628A",
x"7B1E625A",
x"7BA4622F",
x"7C35620B",
x"7CBF61F6",
x"7D2F61F6",
x"7D72620D",
x"7D70623E",
x"7D236284",
x"7C8462D9",
x"7B9E632E",
x"7A826377",
x"794963A7",
x"781163B4",
x"76F76398",
x"760F6356",
x"756062F3",
x"74EA6274",
x"749761E8",
x"744B6152",
x"73E260B8",
x"7334601F",
x"72285F83",
x"70AE5EE0",
x"6ECC5E33",
x"6C9E5D80",
x"6A515CCB",
x"68235C1E",
x"66585B90",
x"65345B35",
x"64EE5B25",
x"65AD5B76",
x"677A5C36",
x"6A4B5D66",
x"6DF85EFE",
x"724560E9",
x"76EB6307",
x"7B9D6534",
x"8016674C",
x"84186930",
x"877C6ACB",
x"8A2E6C13",
x"8C316D10",
x"8D986DD4",
x"8E8E6E78",
x"8F3F6F1C",
x"8FE06FDB",
x"90A470D1",
x"91B4720A",
x"932C738B",
x"951C7548",
x"97817731",
x"9A4A7930",
x"9D577B25",
x"A0837CF7",
x"A3A17E92",
x"A68A7FE6",
x"A91A80F0",
x"AB3B81B2",
x"ACE38235",
x"AE158288",
x"AEE682BD",
x"AF6D82E4",
x"AFC9830C",
x"B019833D",
x"B077837E",
x"B0F583CC",
x"B19E8425",
x"B2708480",
x"B36384D4",
x"B466851E",
x"B5688557",
x"B6598581",
x"B722859C",
x"B7BC85B2",
x"B81F85C8",
x"B84985EA",
x"B841861E",
x"B812866C",
x"B7CC86D3",
x"B7818752",
x"B74587E3",
x"B72C887E",
x"B74A891A",
x"B7A989AC",
x"B8518A31",
x"B93F8AA1",
x"BA648AFD",
x"BBAF8B46",
x"BD048B80",
x"BE408BAE",
x"BF468BD5",
x"BFF78BF6",
x"C03F8C10",
x"C0138C20",
x"BF758C20",
x"BE748C0A",
x"BD268BD6",
x"BBAB8B7E",
x"BA218B00",
x"B8AB8A5A",
x"B7648991",
x"B66088AC",
x"B5A887B9",
x"B54086C3",
x"B52185DC",
x"B53A850D",
x"B57F8464",
x"B5DB83EA",
x"B63A839C",
x"B68B837B",
x"B6C0837B",
x"B6D18392",
x"B6B583B1",
x"B66B83C5",
x"B5F583C3",
x"B557839E",
x"B4978350",
x"B3B682D9",
x"B2BD823D",
x"B1AF8188",
x"B08A80C5",
x"AF4F8000",
x"ADF77F46",
x"AC847EA5",
x"AAEE7E1B",
x"A9397DAD",
x"A7697D59",
x"A5857D14",
x"A39E7CDA",
x"A1C27CA2",
x"A0087C67",
x"9E817C28",
x"9D3D7BE4",
x"9C487B9F",
x"9BA47B5E",
x"9B4B7B28",
x"9B317AFC",
x"9B427ADD",
x"9B697AC4",
x"9B8E7AAA",
x"9B9C7A88",
x"9B887A53",
x"9B497A01",
x"9AE6798F",
x"9A6678FE",
x"99DA7857",
x"995377A3",
x"98E276F4",
x"988A7652",
x"984C75CB",
x"98187561",
x"97D3750C",
x"975974BB",
x"96817457",
x"952273C4",
x"931D72E2",
x"905D719D",
x"8CE36FE5",
x"88C56DBB",
x"842B6B2D",
x"7F51685B",
x"7A7E656F",
x"7600629B",
x"721D6014",
x"6F115E0B",
x"6D075CA2",
x"6C165BF3",
x"6C375C02",
x"6D585CC5",
x"6F515E22",
x"71F05FF6",
x"75026217",
x"7851645C",
x"7BB2669E",
x"7F0368BE",
x"822A6AA6",
x"85186C48",
x"87C96DA3",
x"8A3C6EB5",
x"8C776F8C",
x"8E80702E",
x"905D70AD",
x"92147113",
x"93AA716F",
x"952271CB",
x"967D7233",
x"97BC72AB",
x"98DD7339",
x"99E073DA",
x"9ABF748C",
x"9B7A7546",
x"9C0E75FC",
x"9C7B76A2",
x"9CC27729",
x"9CE77783",
x"9CEE77AA",
x"9CDF7796",
x"9CC17748",
x"9C9A76C6",
x"9C6C7619",
x"9C38754E",
x"9BFD7476",
x"9BB6739F",
x"9B5F72D7",
x"9AF3722A",
x"9A7071A0",
x"99DC7140",
x"993E710C",
x"98A57105",
x"9824712D",
x"97D07182",
x"97BE7200",
x"980172A6",
x"98A9736E",
x"99BE7452",
x"9B3F754D",
x"9D277654",
x"9F647760",
x"A1E17865",
x"A480795D",
x"A71F7A3E",
x"A99A7B05",
x"ABCC7BAA",
x"AD917C29",
x"AED17C81",
x"AF777CAF",
x"AF7B7CB3",
x"AEE67C8F",
x"ADCA7C44",
x"AC4A7BDB",
x"AA927B58",
x"A8CF7AC9",
x"A7337A36",
x"A5E679AD",
x"A504793C",
x"A49978E8",
x"A4A178BC",
x"A50178B6",
x"A59B78D0",
x"A63F7902",
x"A6C0793D",
x"A6F77974",
x"A6C67995",
x"A61E7995",
x"A4FD796E",
x"A373791C",
x"A19778A2",
x"9F857809",
x"9D60775D",
x"9B4276A5",
x"993E75EE",
x"975F753B",
x"95AB7492",
x"942173EE",
x"92B9734D",
x"917072A7",
x"904271F9",
x"8F317143",
x"8E3F7086",
x"8D766FCA",
x"8CDC6F17",
x"8C776E78",
x"8C496DF6",
x"8C4B6D97",
x"8C706D5B",
x"8CA56D3D",
x"8CD26D31",
x"8CDF6D27",
x"8CB26D0F",
x"8C3B6CD8",
x"8B6D6C76",
x"8A4C6BE5",
x"88DD6B23",
x"87356A38",
x"856A6931",
x"839A681D",
x"81D9670E",
x"803E660E",
x"7ED2652A",
x"7D95645F",
x"7C7D63AE",
x"7B74630D",
x"7A5F6272",
x"791D61CF",
x"7793611A",
x"75AD604C",
x"735E5F62",
x"70AD5E5D",
x"6DAB5D48",
x"6A7D5C29",
x"674F5B12",
x"64585A0D",
x"61CB5926",
x"5FDB586A",
x"5EAA57DF",
x"5E4E5788",
x"5ECA5769",
x"600C577E",
x"61EF57C6",
x"6445583D",
x"66D858DF",
x"696D59A6",
x"6BD35A90",
x"6DE55B92",
x"6F875CAE",
x"70B55DD7",
x"71775F0B",
x"71E66041",
x"72206172",
x"724C6297",
x"728D63AA",
x"730064A5",
x"73BA6587",
x"74C4664E",
x"761966FC",
x"77AA6793",
x"79656814",
x"7B2D6886",
x"7CEA68EB",
x"7E846942",
x"7FE9698E",
x"810E69D1",
x"81F36A09",
x"829A6A37",
x"83106A59",
x"835F6A76",
x"83956A8D",
x"83C26AA1",
x"83ED6AB5",
x"841B6ACB",
x"844E6ADC",
x"84806AE9",
x"84AC6AE9",
x"84CE6AD8",
x"84D96AAD",
x"84CB6A66",
x"849E6A03",
x"8456698C",
x"83F7690A",
x"8387688D",
x"83136826",
x"82A467E5",
x"824667D8",
x"82066806",
x"81E9686D",
x"81F66906",
x"822E69BE",
x"828E6A7C",
x"83116B26",
x"83AB6BA3",
x"84526BDE",
x"84F36BCC",
x"85816B69",
x"85ED6ABF",
x"862869E1",
x"862868E9",
x"85EA67F6",
x"85706724",
x"84C2668E",
x"83EC6645",
x"8301664F",
x"821866AA",
x"81436745",
x"809A680D",
x"802A68E6",
x"7FFF69B7",
x"801D6A66",
x"80816AE8",
x"81286B34",
x"82046B4C",
x"83076B3D",
x"84216B13",
x"85466AE3",
x"86656ABD",
x"87736AAB",
x"88656AB5",
x"892E6ADB",
x"89C96B14",
x"8A2F6B55",
x"8A5C6B93",
x"8A4C6BC2",
x"8A036BDB",
x"89866BDC",
x"88DC6BCB",
x"88116BB1",
x"87386B9A",
x"865C6B92",
x"85906BA1",
x"84E26BCF",
x"845A6C17",
x"84036C75",
x"83DA6CD9",
x"83DF6D35",
x"840A6D7D",
x"844E6DA1",
x"84A06D99",
x"84EF6D63",
x"852C6D04",
x"854F6C83",
x"85496BED",
x"85146B4F",
x"84AF6ABA",
x"841B6A34",
x"835A69C5",
x"82796972",
x"817D6935",
x"8074690A",
x"7F6668E8",
x"7E5968C5",
x"7D506894",
x"7C46684E",
x"7B3767E8",
x"7A16675B",
x"78D866A0",
x"777365B5",
x"75E2649B",
x"74256358",
x"724C61F4",
x"706B6081",
x"6EA15F15",
x"6D165DCB",
x"6BF55CBC",
x"6B635C0B",
x"6B875BD0",
x"6C765C1E",
x"6E385D00",
x"70C75E73",
x"74096069",
x"77D962C9",
x"7C06656D",
x"805B682E",
x"84A16AE2",
x"88AD6D66",
x"8C586F9D",
x"8F8E7179",
x"924C72F6",
x"949E7421",
x"969E750D",
x"987075D5",
x"9A3C7699",
x"9C287774",
x"9E56787B",
x"A0D679B9",
x"A3AC7B30",
x"A6CC7CD4",
x"AA157E94",
x"AD598050",
x"B06981EE",
x"B3088350",
x"B509845D",
x"B6478504",
x"B6AF853B",
x"B6438505",
x"B51E8473",
x"B36D8398",
x"B1708291",
x"AF6A817E",
x"ADA2807B",
x"AC577FA2",
x"ABB27F05",
x"ABCC7EB0",
x"ACA37E9F",
x"AE257ED0",
x"B02B7F37",
x"B2827FCA",
x"B4F88080",
x"B75D814F",
x"B98C8235",
x"BB728333",
x"BD0B844F",
x"BE63858D",
x"BF8F86EE",
x"C0AD8876",
x"C1D78A18",
x"C31E8BC9",
x"C48C8D76",
x"C61B8F07",
x"C7B69066",
x"C943917F",
x"CA9D9242",
x"CBA692AA",
x"CC4692B8",
x"CC6D9279",
x"CC1F9200",
x"CB6D9166",
x"CA7590C7",
x"C962903F",
x"C8608FE5",
x"C79B8FC9",
x"C7368FF9",
x"C7449074",
x"C7CD9135",
x"C8C3922E",
x"CA0C9349",
x"CB829472",
x"CCFB958F",
x"CE4B9687",
x"CF56974B",
x"D00297CB",
x"D04D9805",
x"D04397FC",
x"CFFE97BA",
x"CF9F9751",
x"CF5096D6",
x"CF2F965E",
x"CF5795F9",
x"CFD295B1",
x"D098958F",
x"D193958A",
x"D29F959E",
x"D39395BA",
x"D44695CE",
x"D49695CB",
x"D46E95AA",
x"D3CB9565",
x"D2BD94FD",
x"D161947D",
x"CFE093F2",
x"CE6B9368",
x"CD2C92EF",
x"CC469291",
x"CBCE9258",
x"CBCA9244",
x"CC2F924F",
x"CCE29274",
x"CDC092A7",
x"CEA292D9",
x"CF6192FF",
x"CFDB930E",
x"CFF892FC",
x"CFA692C1",
x"CEE49259",
x"CDB091C2",
x"CC1890F9",
x"CA238FFE",
x"C7E08ED5",
x"C5578D7B",
x"C28F8BF3",
x"BF888A3E",
x"BC3C8856",
x"B89E863C",
x"B49E83E6",
x"B025814F",
x"AB227E6E",
x"A5827B3A",
x"9F3B77B2",
x"984F73D5",
x"90CE6FAE",
x"88DD6B52",
x"80AE66DE",
x"78846273",
x"70B15E41",
x"69875A71",
x"63575732",
x"5E6254A5",
x"5ADE52E1",
x"58E251F2",
x"586B51D4",
x"595C5271",
x"5B8553AC",
x"5E9E555D",
x"625F575C",
x"667D5980",
x"6AB75BA4",
x"6ED45DB1",
x"72B15F91",
x"7638613E",
x"796062B4",
x"7C2E63F6",
x"7EA7650D",
x"80D865FD",
x"82C966D1",
x"8481678E",
x"8609683B",
x"875D68DC",
x"88876975",
x"89866A0A",
x"8A626AA1",
x"8B1F6B3A",
x"8BC96BD8",
x"8C676C7A",
x"8CFD6D1D",
x"8D906DBE",
x"8E1E6E55",
x"8EA46EDE",
x"8F1B6F54",
x"8F7C6FB4",
x"8FC16FFE",
x"8FE77031",
x"8FEE7057",
x"8FDC706F",
x"8FB57083",
x"8F847096",
x"8F5270A7",
x"8F2470B9",
x"8EFD70C7",
x"8EDF70CD",
x"8EC570C8",
x"8EAA70B5",
x"8E887094",
x"8E5A7069",
x"8E1C7037",
x"8DCF7008",
x"8D746FE1",
x"8D126FCA",
x"8CAF6FC7",
x"8C536FD7",
x"8C066FFC",
x"8BCB702D",
x"8BA77066",
x"8B9A70A0",
x"8BA470D5",
x"8BC57100",
x"8BFA711F",
x"8C427134",
x"8C9D7140",
x"8D0A714A",
x"8D887154",
x"8E187165",
x"8EB87180",
x"8F6771A7",
x"902471DF",
x"90EA7227",
x"91BC7280",
x"929772E8",
x"937B735F",
x"946A73E1",
x"9564746A",
x"966A74F2",
x"977A7575",
x"988E75EA",
x"99A17646",
x"9AA67681",
x"9B927695",
x"9C55767F",
x"9CE47641",
x"9D3675E0",
x"9D487564",
x"9D1C74DE",
x"9CBC745A",
x"9C3873E8",
x"9BA17393",
x"9B0B7364",
x"9A87735C",
x"9A217378",
x"99E373AF",
x"99CD73F4",
x"99DA743A",
x"9A047476",
x"9A3C74A1",
x"9A7B74BA",
x"9AB874C3",
x"9AF074C8",
x"9B2174D7",
x"9B5274FE",
x"9B88754A",
x"9BCD75C1",
x"9C287664",
x"9C9B772C",
x"9D2B7808",
x"9DD678E7",
x"9E9879AF",
x"9F6D7A50",
x"A0527AB9",
x"A13E7AE4",
x"A2307AD6",
x"A3227A98",
x"A40B7A3A",
x"A4DE79CE",
x"A58A7965",
x"A5F67908",
x"A60078B7",
x"A5857867",
x"A4637806",
x"A2777779",
x"9FAF76A6",
x"9C017574",
x"977873D0",
x"923671B7",
x"8C6A6F31",
x"86586C57",
x"804B6949",
x"7A966638",
x"75806350",
x"714E60C2",
x"6E285EB3",
x"6C285D3D",
x"6B4E5C70",
x"6B825C48",
x"6C9B5CB6",
x"6E685DA5",
x"70AE5EF7",
x"733D608D",
x"75E56249",
x"788A6418",
x"7B1A65E8",
x"7D9467B1",
x"7FFD6970",
x"82636B28",
x"84D26CDB",
x"87556E89",
x"89EA7031",
x"8C8B71CE",
x"8F287352",
x"91A974B4",
x"93F775E4",
x"95FA76D5",
x"979F777E",
x"98DF77DA",
x"99B577E8",
x"9A2977B0",
x"9A48773A",
x"9A1F7696",
x"99BC75CE",
x"992C74F5",
x"98777416",
x"97A2733E",
x"96B17276",
x"95A571C5",
x"94887131",
x"936070BE",
x"923B706B",
x"91287039",
x"903B7024",
x"8F837027",
x"8F0D703B",
x"8EDF7058",
x"8EF97076",
x"8F52708F",
x"8FDD709D",
x"9087709F",
x"913E7094",
x"91F07085",
x"92917075",
x"931A7070",
x"9387707C",
x"93DF70A1",
x"942470E1",
x"945D713D",
x"949271B0",
x"94C37231",
x"94F172BB",
x"95177341",
x"952E73BA",
x"952C7421",
x"950E7472",
x"94D274AD",
x"947774D7",
x"940A74F4",
x"9398750D",
x"9332752A",
x"92F07552",
x"92E3758C",
x"931D75D8",
x"93A87639",
x"948776A9",
x"95B27725",
x"971B77A3",
x"98A9781D",
x"9A427889",
x"9BC878DE",
x"9D217916",
x"9E35792A",
x"9EF6791B",
x"9F5D78E5",
x"9F6A788F",
x"9F257819",
x"9E98778D",
x"9DCF76F2",
x"9CD37650",
x"9BAC75AD",
x"9A5D750D",
x"98E67475",
x"974373E2",
x"95767350",
x"937E72BB",
x"9164721A",
x"8F347169",
x"8D0470A1",
x"8AED6FC3",
x"890D6ED1",
x"87836DD4",
x"86676CDC",
x"85CE6BFA",
x"85C16B42",
x"863B6AC8",
x"87316A9C",
x"88876AC5",
x"8A1D6B44",
x"8BCB6C12",
x"8D676D1A",
x"8ECD6E45",
x"8FE06F79",
x"90877099",
x"90BE7189",
x"90877239",
x"8FF0729A",
x"8F1272AB",
x"8E07726F",
x"8CEC71EC",
x"8BD57131",
x"8ACF7048",
x"89DA6F38",
x"88ED6E08",
x"87EF6CB8",
x"86C36B47",
x"854B69B0",
x"836667F3",
x"81046613",
x"7E1E6414",
x"7ABE6204",
x"76FD5FF4",
x"73075DF8",
x"6F0C5C22",
x"6B445A87",
x"67E25935",
x"65135833",
x"62F65787",
x"619A572B",
x"61025717",
x"611B5740",
x"61D2579B",
x"6305581C",
x"649458BC",
x"66625975",
x"68585A43",
x"6A635B24",
x"6C785C14",
x"6E915D12",
x"70AA5E1A",
x"72C15F22",
x"74D56024",
x"76E26117",
x"78E361F6",
x"7AD262BB",
x"7CAB6368",
x"7E6D6403",
x"80176493",
x"81AE6523",
x"833865C1",
x"84C16677",
x"8652674E",
x"87F46846",
x"89AE6962",
x"8B7D6A96",
x"8D5B6BD7",
x"8F3E6D1A",
x"91146E4F",
x"92C96F6C",
x"94487064",
x"957D7133",
x"965C71D7",
x"96DA724D",
x"96FB729A",
x"96C872C3",
x"965072CA",
x"95AB72B6",
x"94F4728A",
x"94497250",
x"93C8720D",
x"938771CA",
x"939E7195",
x"941B7178",
x"95037183",
x"965671C3",
x"980D723E",
x"9A1472FB",
x"9C5973F6",
x"9EBF7527",
x"A129767E",
x"A37877E5",
x"A58F7947",
x"A7567A8C",
x"A8BD7BA0",
x"A9BB7C77",
x"AA4D7D09",
x"AA7E7D59",
x"AA5D7D6B",
x"AA007D51",
x"A97D7D18",
x"A8E97CD0",
x"A8597C88",
x"A7DC7C49",
x"A77A7C1B",
x"A7397BFC",
x"A7197BEF",
x"A7197BEE",
x"A7367BF7",
x"A76A7C05",
x"A7B27C19",
x"A80D7C30",
x"A8757C49",
x"A8E77C64",
x"A95D7C7E",
x"A9CF7C95",
x"AA367CA3",
x"AA8B7CA5",
x"AACA7C96",
x"AAEE7C78",
x"AAFB7C4A",
x"AAF37C11",
x"AAD97BD6",
x"AAB67B9F",
x"AA8A7B77",
x"AA537B61",
x"AA0C7B60",
x"A9AE7B72",
x"A9297B8F",
x"A8737BAD",
x"A7857BBF",
x"A65E7BB9",
x"A5077B93",
x"A3907B4D",
x"A2127AE5",
x"A0AB7A68",
x"9F7779E3",
x"9E8D7962",
x"9DF878F5",
x"9DB978A3",
x"9DC27871",
x"9DF7785A",
x"9E357854",
x"9E57784D",
x"9E397836",
x"9DC077FC",
x"9CE17796",
x"9B9B76FB",
x"99FE7630",
x"9824753D",
x"96297431",
x"942C731D",
x"92437212",
x"90767116",
x"8EC17031",
x"8D106F59",
x"8B456E86",
x"893E6DA4",
x"86DD6CA3",
x"840A6B70",
x"80C26A07",
x"7D13686C",
x"792166AB",
x"752864E0",
x"716D632F",
x"6E3B61BB",
x"6BDB60A9",
x"6A876018",
x"6A626015",
x"6B7860A4",
x"6DB561B5",
x"70F0632F",
x"74E964ED",
x"795566C6",
x"7DE96894",
x"82606A37",
x"86846B9A",
x"8A326CB7",
x"8D5C6D90",
x"90046E38",
x"92406ECA",
x"942C6F61",
x"95E77017",
x"97907106",
x"9940723B",
x"9B0A73B9",
x"9CF7757B",
x"9F0A7771",
x"A13F7988",
x"A3927BA6",
x"A5F77DB0",
x"A8637F91",
x"AAC58133",
x"AD0B828E",
x"AF1F8397",
x"B0EE844D",
x"B26184B9",
x"B36384E1",
x"B3E884D0",
x"B3F08494",
x"B37E8433",
x"B2A883B8",
x"B1878326",
x"B0408282",
x"AEF581CF",
x"ADC9810C",
x"ACD3803D",
x"AC1B7F67",
x"ABA37E91",
x"AB5D7DC1",
x"AB317D06",
x"AB047C6A",
x"AABB7BF5",
x"AA427BB3",
x"A98E7BA2",
x"A89F7BC0",
x"A77E7C04",
x"A63C7C5E",
x"A4EE7CBF",
x"A3AB7D0E",
x"A2827D3C",
x"A1817D3C",
x"A0AF7D04",
x"A00A7C96",
x"9F8E7BFB",
x"9F357B3E",
x"9EF77A78",
x"9ED079BC",
x"9EBF7920",
x"9EC678B9",
x"9EE77890",
x"9F2478AC",
x"9F80790B",
x"9FF979A0",
x"A08D7A5E",
x"A1367B30",
x"A1F17C01",
x"A2B57CBD",
x"A3807D54",
x"A4497DBC",
x"A5117DEE",
x"A5D27DEE",
x"A6877DC0",
x"A72B7D6E",
x"A7B67D02",
x"A81E7C89",
x"A8577C0C",
x"A8567B95",
x"A8157B29",
x"A78F7ACA",
x"A6C97A79",
x"A5CA7A37",
x"A4A17A01",
x"A36179D3",
x"A21E79AD",
x"A0EA798C",
x"9FD2796D",
x"9EE07950",
x"9E177932",
x"9D737915",
x"9CED78F9",
x"9C7D78E0",
x"9C1B78CD",
x"9BC278C4",
x"9B7478CD",
x"9B3578E8",
x"9B0D791C",
x"9B07796A",
x"9B2B79D0",
x"9B807A47",
x"9C047AC9",
x"9CAF7B46",
x"9D747BB4",
x"9E3F7C02",
x"9EFA7C25",
x"9F8E7C13",
x"9FEC7BCD",
x"A0087B56",
x"9FE37AB7",
x"9F807A01",
x"9EEA7941",
x"9E317889",
x"9D5A77E1",
x"9C6E774A",
x"9B6376BE",
x"9A29762D",
x"98A4757E",
x"96AF7495",
x"94287357",
x"90F071AD",
x"8CF46F8C",
x"88376CF6",
x"82D269FF",
x"7CF666C6",
x"76ED637C",
x"710C6050",
x"6BAE5D7D",
x"672A5B2F",
x"63C7598B",
x"61B458A6",
x"61005882",
x"619C590F",
x"635C5A2C",
x"65FC5BB3",
x"692B5D73",
x"6C965F3F",
x"6FEF60F0",
x"72F7626C",
x"7587639F",
x"778C648A",
x"7907652F",
x"7A0D65A1",
x"7ABB65F2",
x"7B346635",
x"7B97667A",
x"7C0066CF",
x"7C7F673A",
x"7D1A67B8",
x"7DD06848",
x"7E9B68DF",
x"7F6F6975",
x"804269FF",
x"810A6A75",
x"81C26AD1",
x"82666B11",
x"82F46B37",
x"836F6B47",
x"83D26B44",
x"841D6B37",
x"84496B27",
x"84526B1C",
x"842F6B19",
x"83DF6B21",
x"835A6B37",
x"82A86B55",
x"81CB6B78",
x"80D16B96",
x"7FC86BA8",
x"7EC56BA7",
x"7DD66B8A",
x"7D0D6B4F",
x"7C736AF6",
x"7C0D6A80",
x"7BD869F5",
x"7BCC695F",
x"7BE268C8",
x"7C0A683F",
x"7C3967CB",
x"7C696775",
x"7C93673E",
x"7CB76727",
x"7CD96727",
x"7CFD6735",
x"7D286746",
x"7D5F674F",
x"7D9E6744",
x"7DE5671E",
x"7E2D66DE",
x"7E6F6686",
x"7EA5661E",
x"7ECF65B8",
x"7EF0655F",
x"7F116527",
x"7F3E651B",
x"7F866549",
x"7FFA65B4",
x"80A56659",
x"818B6732",
x"82AD6831",
x"83FD6941",
x"856A6A4E",
x"86DF6B41",
x"88416C06",
x"897A6C8D",
x"8A7C6CCD",
x"8B396CC4",
x"8BB46C78",
x"8BF16BF6",
x"8C006B52",
x"8BEC6AA6",
x"8BC56A06",
x"8B9A698C",
x"8B6F6945",
x"8B48693C",
x"8B216973",
x"8AF369E1",
x"8AB56A76",
x"8A626B21",
x"89F46BCA",
x"896C6C5F",
x"88D06CD1",
x"88286D19",
x"87836D37",
x"86ED6D31",
x"86716D14",
x"861D6CEE",
x"85F06CCB",
x"85E96CB7",
x"85FE6CB4",
x"86256CBF",
x"86496CD2",
x"86596CE1",
x"86456CD9",
x"85FE6CB4",
x"85816C68",
x"84CE6BF5",
x"83EF6B61",
x"82F76ABA",
x"82006A11",
x"8122697A",
x"80776907",
x"801368C1",
x"7FFC68AD",
x"802D68C2",
x"808D68F3",
x"80FA6928",
x"81416944",
x"81286927",
x"807668B5",
x"7EFA67DE",
x"7C916690",
x"793164CE",
x"74E362A2",
x"6FD46022",
x"6A3F5D6A",
x"64795AA1",
x"5ED957E9",
x"59BE5566",
x"55785339",
x"52445178",
x"504A5035",
x"4F944F75",
x"50184F39",
x"51AB4F77",
x"5419501C",
x"571E5116",
x"5A78524A",
x"5DE253A2",
x"61275501",
x"641A5654",
x"66A0578A",
x"68A85894",
x"6A37596E",
x"6B535A18",
x"6C115A9B",
x"6C895B00",
x"6CD45B56",
x"6D0C5BAB",
x"6D445C0D",
x"6D8C5C87",
x"6DEE5D1A",
x"6E695DC5",
x"6EFC5E81",
x"6F995F43",
x"70375FFC",
x"70C5609B",
x"713A611A",
x"718C6170",
x"71B7619B",
x"71C161A2",
x"71B0618D",
x"718C6169",
x"71636141",
x"713E611F",
x"7124610B",
x"71166103",
x"71136100",
x"711460FC",
x"711460E9",
x"710C60BE",
x"70F66076",
x"70D2600D",
x"70A65F8D",
x"70775F00",
x"70555E78",
x"70485E0B",
x"70595DCD",
x"70935DCC",
x"70F05E11",
x"71705E9E",
x"72065F67",
x"72A3605F",
x"7334616C",
x"73AA6277",
x"73F86366",
x"74166424",
x"73FF64A4",
x"73BA64DE",
x"734F64D2",
x"72CC648B",
x"7242641A",
x"71BF638E",
x"715262FA",
x"71046273",
x"70DC6203",
x"70DB61B4",
x"70FC618A",
x"713B6183",
x"7191619B",
x"71F761C8",
x"72686204",
x"72DC6243",
x"73526281",
x"73C762B9",
x"743962EA",
x"74A86315",
x"7511633C",
x"75706362",
x"75C26387",
x"760063AA",
x"762863C8",
x"763463DC",
x"762463DF",
x"75F663CB",
x"75AE639B",
x"75516350",
x"74E262EF",
x"74696280",
x"73F06211",
x"737A61B2",
x"73116173",
x"72B86163",
x"7275618A",
x"724B61E8",
x"723E6274",
x"724C6324",
x"727963E0",
x"72BF6494",
x"731E6528",
x"738E658D",
x"740A65B4",
x"7486659E",
x"74FA6552",
x"755B64DC",
x"75A1644F",
x"75C663C2",
x"75C86345",
x"75A562EA",
x"756362B7",
x"750762AD",
x"749762C2",
x"741E62ED",
x"739E631B",
x"731D633C",
x"7297633E",
x"720A6313",
x"716B62B1",
x"70B06215",
x"6FCB6141",
x"6EB26035",
x"6D5B5EFC",
x"6BC15D9C",
x"69E35C22",
x"67CB5A98",
x"6583590A",
x"631D577F",
x"60B05609",
x"5E5754AF",
x"5C2A537E",
x"5A44527F",
x"58BE51BD",
x"57AA513D",
x"57165104",
x"5709510F",
x"577F5160",
x"587051EA",
x"59CA52A5",
x"5B725385",
x"5D4B547A",
x"5F35557A",
x"61115675",
x"62C45767",
x"64385846",
x"65625911",
x"663F59C6",
x"66DB5A67",
x"67455AFA",
x"67975B7E",
x"67EC5BF8",
x"685C5C6A",
x"68FB5CD6",
x"69D15D3C",
x"6ADE5D9C",
x"6C175DF7",
x"6D685E4C",
x"6EB25E9F",
x"6FDE5EF0",
x"70CB5F41",
x"71685F92",
x"71A75FE6",
x"718A6038",
x"71196086",
x"706560CB",
x"6F8A6101",
x"6EA36124",
x"6DC9612E",
x"6D14611E",
x"6C9360F0",
x"6C4F60A9",
x"6C49604F",
x"6C7A5FE3",
x"6CDB5F72",
x"6D585EFE",
x"6DE55E8E",
x"6E705E25",
x"6EEB5DC5",
x"6F4B5D6C",
x"6F865D18",
x"6F975CCB",
x"6F7F5C81",
x"6F415C3C",
x"6EE35C00",
x"6E755BD3",
x"6E025BBC",
x"6D9A5BC3",
x"6D4F5BEE",
x"6D305C40",
x"6D475CB9",
x"6D9A5D53",
x"6E2E5E04",
x"6EFA5EC1",
x"6FF55F77",
x"710E601A",
x"7232609B",
x"734B60F0",
x"74476115",
x"7511610A",
x"75A060D5",
x"75EA607D",
x"75F26011",
x"75BC5F9E",
x"75545F2C",
x"74C75ECB",
x"74275E7E",
x"73845E4B",
x"72EF5E31",
x"72725E32",
x"72115E4C",
x"71D15E7A",
x"71AE5EB9",
x"71A45F0A",
x"71AA5F66",
x"71B85FC9",
x"71C86031",
x"71D56097",
x"71DB60F4",
x"71D96143",
x"71D3617D",
x"71CB619D",
x"71C461A1",
x"71BF618A",
x"71BE615C",
x"71BF611D",
x"71BF60D5",
x"71B8608D",
x"71A7604B",
x"71846015",
x"714E5FF0",
x"71035FD8",
x"70A35FCC",
x"70305FC9",
x"6FAE5FC6",
x"6F245FC3",
x"6E965FBB",
x"6E095FAB",
x"6D825F98",
x"6D045F81",
x"6C935F69",
x"6C315F50",
x"6BDF5F39",
x"6B9D5F21",
x"6B6C5F03",
x"6B495EDC",
x"6B305EA7",
x"6B175E5F",
x"6AF65E00",
x"6AC15D8B",
x"6A6B5D04",
x"69EC5C70",
x"693B5BD5",
x"685C5B3F",
x"67565AB9",
x"663D5A4D",
x"65285A05",
x"643B59EA",
x"639A5A04",
x"63665A53",
x"63BD5ADA",
x"64AE5B97",
x"663E5C84",
x"68605D9E",
x"6B005EDA",
x"6DF86033",
x"7120619F",
x"74536317",
x"776D6495",
x"7A596616",
x"7D0A6796",
x"7F846913",
x"81D36A8D",
x"840E6C04",
x"864C6D79",
x"88A76EE8",
x"8B2C704F",
x"8DE671AF",
x"90D57302",
x"93EA7447",
x"9718757B",
x"9A46769C",
x"9D5C77A9",
x"A04578A3",
x"A2EB798C",
x"A5437A63",
x"A7437B29",
x"A8E77BE1",
x"AA307C89",
x"AB227D20",
x"ABC27DA3",
x"AC177E11",
x"AC2B7E64",
x"AC087E9C",
x"ABB97EB3",
x"AB477EAD",
x"AAC27E88",
x"AA2E7E47",
x"A9957DEF",
x"A8FB7D85",
x"A8637D0E",
x"A7C97C8F",
x"A72B7C0E",
x"A6847B8C",
x"A5D07B0E",
x"A5127A96",
x"A44A7A29",
x"A38779C6",
x"A2D37972",
x"A2467933",
x"A1F4790C",
x"A1F07901",
x"A2487915",
x"A302794A",
x"A418799B",
x"A5777A05",
x"A7037A81",
x"A8947B01",
x"AA027B7E",
x"AB297BEA",
x"ABEA7C3D",
x"AC327C74",
x"AC047C8B",
x"AB717C86",
x"AA9B7C6E",
x"A9B07C4A",
x"A8E37C29",
x"A8647C15",
x"A85C7C19",
x"A8DF7C3A",
x"A9F37C7C",
x"AB847CDB",
x"AD707D51",
x"AF8A7DD1",
x"B1947E51",
x"B35A7EC3",
x"B4AB7F18",
x"B5617F49",
x"B56D7F4C",
x"B4CA7F20",
x"B3887EC9",
x"B1C57E4A",
x"AFA57DB0",
x"AD4F7D05",
x"AAEA7C59",
x"A8947BB6",
x"A6647B28",
x"A4677AB6",
x"A2A27A64",
x"A1127A32",
x"9FAE7A18",
x"9E6D7A12",
x"9D497A16",
x"9C3D7A1D",
x"9B4F7A1D",
x"9A807A15",
x"99DC79FC",
x"996A79D7",
x"993479A6",
x"9939796D",
x"9976792D",
x"99DF78ED",
x"9A6078AA",
x"9AE37865",
x"9B49781C",
x"9B7D77CD",
x"9B667771",
x"9AF97705",
x"9A317688",
x"991775F8",
x"97BE7555",
x"963974A3",
x"94AA73E4",
x"9325731F",
x"91C57257",
x"90937190",
x"8F9170CB",
x"8EB27009",
x"8DE06F45",
x"8CFA6E78",
x"8BDC6D99",
x"8A606C9E",
x"88676B82",
x"85DC6A37",
x"82B868BE",
x"7F046714",
x"7ADE6542",
x"766F6352",
x"71EF6156",
x"6D9E5F63",
x"69BC5D90",
x"66845BF3",
x"64235AA4",
x"62B659AF",
x"62455924",
x"62C75900",
x"641A5943",
x"661459E3",
x"68805ACF",
x"6B285BF8",
x"6DD85D4B",
x"70685EB7",
x"72BD6031",
x"74CE61AB",
x"769B6323",
x"78346493",
x"79AA65F9",
x"7B146752",
x"7C83689B",
x"7E0069D1",
x"7F916AE9",
x"812D6BDC",
x"82C86CA4",
x"844F6D38",
x"85B26D99",
x"86E36DC5",
x"87D66DC4",
x"888B6D9E",
x"89066D63",
x"894F6D1D",
x"89736CD8",
x"897D6C9C",
x"897A6C6C",
x"89706C47",
x"89636C2A",
x"89526C0D",
x"89396BEB",
x"89146BB8",
x"88DC6B76",
x"888B6B23",
x"88206ABF",
x"87986A54",
x"86F669E2",
x"863B6972",
x"856A6909",
x"848968AA",
x"839D6856",
x"82AE6810",
x"81C667DB",
x"80F267B7",
x"803C67A8",
x"7FB267B5",
x"7F5D67E3",
x"7F456835",
x"7F6968AB",
x"7FC26944",
x"804169F5",
x"80D16AB1",
x"81596B68",
x"81BE6C06",
x"81E96C78",
x"81CB6CB3",
x"815F6CAD",
x"80AA6C66",
x"7FC16BE6",
x"7EBC6B3F",
x"7DBF6A82",
x"7CED69C4",
x"7C636919",
x"7C376891",
x"7C706838",
x"7D09680E",
x"7DEF6810",
x"7F066832",
x"80276869",
x"812E68A4",
x"81F968D6",
x"826F68F5",
x"828168F7",
x"822F68D9",
x"8186689E",
x"80986849",
x"7F8467E2",
x"7E676770",
x"7D5E66FA",
x"7C7C6689",
x"7BCE6621",
x"7B5B65C4",
x"7B1B6575",
x"7B066531",
x"7B0764F7",
x"7B1164C4",
x"7B106491",
x"7AF96460",
x"7AC4642A",
x"7A6D63F0",
x"79F763B4",
x"79666376",
x"78C4633C",
x"7817630A",
x"776962E4",
x"76BF62D0",
x"761E62CC",
x"758A62D5",
x"750362E8",
x"748762FC",
x"7419630A",
x"73B16307",
x"735262F0",
x"72F962C1",
x"72A76277",
x"725B621D",
x"721861B7",
x"71E16150",
x"71B860F3",
x"719E60A9",
x"71936074",
x"71906056",
x"718C6049",
x"717A6042",
x"71486037",
x"70E5601A",
x"703C5FDD",
x"6F445F7D",
x"6DF35EF4",
x"6C4F5E46",
x"6A665D7A",
x"68525C9C",
x"66315BB9",
x"642B5AE1",
x"62665A21",
x"61035982",
x"601A590C",
x"5FB758C3",
x"5FD858A5",
x"606F58AF",
x"616558DD",
x"62995928",
x"63EB598A",
x"653E59FB",
x"66785A77",
x"678A5AF7",
x"686C5B74",
x"69205BEC",
x"69A85C55",
x"6A105CAE",
x"6A615CF4",
x"6AA05D24",
x"6AD55D3F",
x"6B025D48",
x"6B275D46",
x"6B475D41",
x"6B655D42",
x"6B865D55",
x"6BB25D86",
x"6BF65DDA",
x"6C595E5A",
x"6CE95F06",
x"6DA95FD9",
x"6E9A60CC",
x"6FB561D2",
x"70F062DA",
x"723863D5",
x"737864B1",
x"74966560",
x"758165D9",
x"762D6616",
x"768F661A",
x"76A865E9",
x"7684658D",
x"76326513",
x"75C66489",
x"755B63F9",
x"7500636F",
x"74CE62F4",
x"74CE6290",
x"75096245",
x"757F621A",
x"762A6210",
x"76FF622B",
x"77F26270",
x"78F262E2",
x"79F26381",
x"7AE5644E",
x"7BBF6542",
x"7C776653",
x"7D0B6775",
x"7D776891",
x"7DBE6994",
x"7DE26A68",
x"7DE86AFC",
x"7DD86B44",
x"7DB86B3B",
x"7D906AE6",
x"7D626A52",
x"7D316994",
x"7D0068C4",
x"7CCE67FA",
x"7C97674C",
x"7C5966CB",
x"7C13667A",
x"7BC1665E",
x"7B656669",
x"7B046690",
x"7AA166C2",
x"7A4466F0",
x"79F36710",
x"79B56719",
x"7990670D",
x"798366EF",
x"798E66C8",
x"79AA66A1",
x"79CE667F",
x"79EF6665",
x"7A026650",
x"79FC663E",
x"79D66623",
x"798D65F5",
x"792165A8",
x"7896653A",
x"77F364A5",
x"774263F3",
x"768D632D",
x"75DC625F",
x"753A619B",
x"74AA60F2",
x"742F606E",
x"73CE601B",
x"73825FF7",
x"73486001",
x"7321602F",
x"73076074",
x"72F960C1",
x"72F56106",
x"72F96138",
x"7302614F",
x"730E6145",
x"731D611D",
x"732760DA",
x"732A6087",
x"7321602D",
x"73045FD6",
x"72D15F8E",
x"72805F59",
x"720E5F3B",
x"717A5F31",
x"70C25F37",
x"6FE65F43",
x"6EEC5F4F",
x"6DD85F4F",
x"6CB45F3B",
x"6B875F0D",
x"6A5C5EC3",
x"693B5E5D",
x"682D5DDF",
x"67385D4C",
x"66655CAE",
x"65B75C08",
x"65335B67",
x"64E25AD0",
x"64CD5A50",
x"650259F1",
x"658F59BF",
x"668459C9",
x"67F55A1E",
x"69EC5AC9",
x"6C6F5BD6",
x"6F795D46",
x"72FA5F18",
x"76D4613C",
x"7ADC639E",
x"7EE56620",
x"82B9689E",
x"862C6AF9",
x"89176D0D",
x"8B656EC4",
x"8D107013",
x"8E2870F8",
x"8EC97180",
x"8F1D71C3",
x"8F4B71DA",
x"8F7D71E5",
x"8FD57202",
x"90647241",
x"912E72AF",
x"92287348",
x"933B7403",
x"944D74CE",
x"9541758D",
x"95FD762D",
x"96747695",
x"96A476B7",
x"96917690",
x"964D7620",
x"95EE7572",
x"95887499",
x"953273A6",
x"94F672B0",
x"94D771CA",
x"94D67100",
x"94E37061",
x"94F16FEF",
x"94EF6FAE",
x"94CC6F9A",
x"94816FB0",
x"940B6FE8",
x"9371703B",
x"92C070A6",
x"9207711D",
x"9158719C",
x"90C5721A",
x"9058728C",
x"901572EB",
x"8FF97329",
x"8FF4733B",
x"8FF6731A",
x"8FE972BE",
x"8FB37224",
x"8F48714F",
x"8E9A7048",
x"8DA86F1A",
x"8C7B6DD8",
x"8B256C96",
x"89BC6B66",
x"885D6A5C",
x"87226986",
x"862068EC",
x"85656893",
x"84F66876",
x"84CF688D",
x"84E068CE",
x"85176928",
x"855F6993",
x"85A06A02",
x"85C66A6B",
x"85C86AC9",
x"859E6B1D",
x"854B6B63",
x"84D66B9E",
x"844B6BCE",
x"83BC6BF2",
x"83376C09",
x"82CC6C13",
x"82876C0F",
x"826F6BFA",
x"82896BD7",
x"82D36BA7",
x"834E6B70",
x"83F06B3A",
x"84B26B0C",
x"858B6AEC",
x"86706AE3",
x"87566AF3",
x"88346B1E",
x"88FD6B62",
x"89A96BB7",
x"8A356C16",
x"8A9B6C78",
x"8AD86CD1",
x"8AEC6D1C",
x"8ADA6D4F",
x"8AA76D6B",
x"8A556D6E",
x"89E96D59",
x"896A6D33",
x"88DA6CFD",
x"883F6CBE",
x"87976C7A",
x"86E56C33",
x"862B6BE9",
x"85696B9D",
x"84A26B4E",
x"83DD6AF7",
x"831E6A9C",
x"826F6A3A",
x"81D569D5",
x"81586972",
x"80FA6917",
x"80B968C8",
x"808C6889",
x"805F6856",
x"8016682D",
x"7F8D67FD",
x"7EA067B7",
x"7D256742",
x"7AFC6687",
x"780C656C",
x"744E63E2",
x"6FCE61DD",
x"6AAB5F62",
x"651C5C80",
x"5F645955",
x"59D25608",
x"54B752CC",
x"505F4FD3",
x"4D054D4B",
x"4AD14B5E",
x"49D14A26",
x"49FC49AD",
x"4B3049EF",
x"4D384AD8",
x"4FD54C44",
x"52C54E0E",
x"55C85008",
x"58AE520C",
x"5B5153F7",
x"5D9D55AF",
x"5F925729",
x"61355860",
x"629C5959",
x"63DB5A1E",
x"65065ABB",
x"662D5B3B",
x"67595BA9",
x"688C5C0A",
x"69C05C60",
x"6AEB5CAE",
x"6C025CEE",
x"6CF85D24",
x"6DC75D4C",
x"6E6A5D6A",
x"6EE25D84",
x"6F325D9F",
x"6F655DC3",
x"6F835DF4",
x"6F965E38",
x"6FA75E8D",
x"6FBB5EF0",
x"6FD65F5A",
x"6FF75FC2",
x"7019601D",
x"70346060",
x"703F6084",
x"70306084",
x"6FFF605F",
x"6FA16015",
x"6F145FAE",
x"6E555F31",
x"6D695EA4",
x"6C565E10",
x"6B2B5D7B",
x"69F55CEC",
x"68C55C64",
x"67B05BE7",
x"66C25B76",
x"660C5B11",
x"65945ABB",
x"655E5A71",
x"65655A39",
x"65A15A12",
x"660459FE",
x"667C59FA",
x"66F55A02",
x"675F5A17",
x"67AD5A32",
x"67D45A52",
x"67D45A73",
x"67B05A95",
x"67735AB9",
x"67305AE4",
x"66F65B18",
x"66DB5B5A",
x"66EE5BAF",
x"67385C17",
x"67BF5C90",
x"687F5D15",
x"69695DA4",
x"6A6D5E33",
x"6B755EBC",
x"6C665F37",
x"6D2B5F9F",
x"6DB35FF2",
x"6DF0602D",
x"6DE36052",
x"6D916062",
x"6D0C605F",
x"6C65604C",
x"6BB7602E",
x"6B1C6007",
x"6AAB5FDF",
x"6A795FB9",
x"6A905F9E",
x"6AF65F91",
x"6BA45F9A",
x"6C905FB9",
x"6DA55FED",
x"6ECF602F",
x"6FF36079",
x"70F960BC",
x"71CC60EC",
x"725F60FC",
x"72A760E4",
x"72A360A4",
x"725D603C",
x"71E25FB9",
x"71455F2B",
x"709D5EA4",
x"6FFF5E36",
x"6F7D5DF3",
x"6F255DDF",
x"6EFD5DFD",
x"6F045E45",
x"6F305EA7",
x"6F735F0E",
x"6FBC5F67",
x"6FFA5F9D",
x"701D5FA1",
x"70195F6E",
x"6FE85F07",
x"6F895E74",
x"6F025DC6",
x"6E595D0E",
x"6D945C5F",
x"6CBA5BC5",
x"6BC85B47",
x"6ABF5AE7",
x"69995A9C",
x"684B5A5A",
x"66CE5A0E",
x"651E59A8",
x"633B591A",
x"612D585C",
x"5F04576B",
x"5CD95651",
x"5AC7551E",
x"58EC53E8",
x"576952C9",
x"565551DB",
x"55C45139",
x"55C050F1",
x"56485111",
x"57575198",
x"58D8527F",
x"5AB753B6",
x"5CDB5526",
x"5F2756B6",
x"6180584D",
x"63D259D0",
x"66075B2F",
x"68105C5F",
x"69E35D57",
x"6B7D5E1C",
x"6CDF5EB3",
x"6E0C5F29",
x"6F0C5F87",
x"6FED5FD9",
x"70BC6029",
x"71876080",
x"725660DF",
x"73356148",
x"742561BB",
x"75256235",
x"763262B4",
x"77416337",
x"784563B9",
x"7935643C",
x"7A0A64BB",
x"7ABD6532",
x"7B4B65A0",
x"7BB965FD",
x"7C0E6644",
x"7C53666D",
x"7C8D6677",
x"7CC4665E",
x"7CF76624",
x"7D2865CC",
x"7D4C6563",
x"7D5C64F4",
x"7D4E648B",
x"7D196438",
x"7CB86407",
x"7C2D63FF",
x"7B806425",
x"7AC16477",
x"7A0364EF",
x"795C6580",
x"78E6661D",
x"78B166B5",
x"78CB673C",
x"793767A7",
x"79F267EC",
x"7AEC680A",
x"7C136804",
x"7D4F67E2",
x"7E8967AE",
x"7FAA6773",
x"80A46741",
x"8170671E",
x"820D6716",
x"8281672D",
x"82DE675F",
x"832B67AB",
x"837D6809",
x"83DA686C",
x"844C68CB",
x"84D06919",
x"8560694C",
x"85F46965",
x"867E695E",
x"86F1693F",
x"87426911",
x"876D68E1",
x"876F68BC",
x"874968B4",
x"870668D4",
x"86AC6920",
x"8646699D",
x"85DD6A45",
x"85766B0C",
x"85116BE1",
x"84AF6CAE",
x"84496D5E",
x"83DC6DDE",
x"835F6E1D",
x"82D06E13",
x"822D6DBD",
x"81766D20",
x"80B46C4A",
x"7FEF6B4B",
x"7F316A3B",
x"7E87692E",
x"7DFF6838",
x"7D9D676D",
x"7D6866D8",
x"7D60667D",
x"7D81665F",
x"7DC46677",
x"7E1866BB",
x"7E726720",
x"7EC16794",
x"7EF5680A",
x"7F046876",
x"7EE668CB",
x"7E976901",
x"7E176916",
x"7D696904",
x"7C9768D1",
x"7BA8687D",
x"7AA4680E",
x"79906787",
x"786C66EC",
x"7737663E",
x"75E86579",
x"7476649D",
x"72D563A7",
x"70FC6293",
x"6EE6615F",
x"6C976010",
x"6A1D5EAB",
x"678D5D3D",
x"65095BD7",
x"62BA5A8B",
x"60CC5973",
x"5F6B58A2",
x"5EBE582E",
x"5EE45828",
x"5FEB589A",
x"61D55988",
x"64945AED",
x"680D5CC1",
x"6C195EEE",
x"70866160",
x"752463FA",
x"79C466A3",
x"7E37693C",
x"825C6BAD",
x"86166DDE",
x"89526FC1",
x"8C0B714D",
x"8E43727F",
x"9003735E",
x"915973F6",
x"925A745B",
x"931F749F",
x"93C074D4",
x"9453750F",
x"94EC7558",
x"959775B6",
x"965D7626",
x"974076A0",
x"98397718",
x"993F777E",
x"9A4077C6",
x"9B3177E5",
x"9C0177DD",
x"9CAB77AC",
x"9D277761",
x"9D787709",
x"9DA476B6",
x"9DB27677",
x"9DAE7658",
x"9D9C7662",
x"9D84768F",
x"9D6976D8",
x"9D48772F",
x"9D1C777C",
x"9CE377AF",
x"9C9877B6",
x"9C397786",
x"9BC8771D",
x"9B48767C",
x"9ABE75B4",
x"9A3274D5",
x"99AC73F8",
x"99317334",
x"98C0729F",
x"985C7248",
x"98007239",
x"97A77270",
x"974B72E8",
x"96E7738F",
x"9678744D",
x"95FC750B",
x"957075B0",
x"94D57626",
x"942F7660",
x"93837651",
x"92D375FF",
x"9227756E",
x"918074AC",
x"90E673CA",
x"905A72DB",
x"8FE271EE",
x"8F7D7112",
x"8F2C704E",
x"8EED6FA9",
x"8EBC6F21",
x"8E946EB8",
x"8E6D6E6B",
x"8E456E35",
x"8E146E1C",
x"8DDB6E1A",
x"8D986E35",
x"8D4F6E6C",
x"8D016EBB",
x"8CB86F23",
x"8C736F97",
x"8C35700F",
x"8BFD707E",
x"8BCB70D7",
x"8B95710F",
x"8B5D7120",
x"8B1B7108",
x"8AD370C8",
x"8A87706B",
x"8A3F6FFE",
x"8A066F8F",
x"89E46F2E",
x"89E66EE6",
x"8A0E6EC1",
x"8A5D6EC5",
x"8ACC6EF0",
x"8B4E6F41",
x"8BD06FAE",
x"8C43702E",
x"8C9370B7",
x"8CB1713A",
x"8C9871AD",
x"8C487205",
x"8BC67237",
x"8B217240",
x"8A67721A",
x"89AF71C7",
x"8908714E",
x"888370BA",
x"882B701A",
x"88086F82",
x"881E6F05",
x"886A6EB4",
x"88E36E9C",
x"897C6EC1",
x"8A1F6F1C",
x"8AB66F9C",
x"8B1E7026",
x"8B357097",
x"8AD370CA",
x"89D97097",
x"882A6FE2",
x"85B56E97",
x"827E6CB5",
x"7E9A6A49",
x"7A316776",
x"75796466",
x"70BB6152",
x"6C3E5E70",
x"684B5BF8",
x"651E5A17",
x"62E358E4",
x"61B4586E",
x"619058AE",
x"6263598B",
x"640D5AE7",
x"665C5C9A",
x"69205E77",
x"6C26605C",
x"6F446228",
x"725663C5",
x"75446528",
x"77F9664B",
x"7A6D6730",
x"7C9567D9",
x"7E6C684E",
x"7FEC6894",
x"811168B0",
x"81D968A4",
x"82486877",
x"825F682D",
x"822E67CF",
x"81C36768",
x"81346706",
x"809766B8",
x"7FFF668D",
x"7F7F6690",
x"7F2266C8",
x"7EEF6737",
x"7EE367D8",
x"7EF5689B",
x"7F1B6973",
x"7F466A47",
x"7F6C6B00",
x"7F806B8C",
x"7F7F6BD8",
x"7F676BDE",
x"7F3C6B99",
x"7F036B10",
x"7EC86A4F",
x"7E906969",
x"7E676875",
x"7E536787",
x"7E5866B8",
x"7E766618",
x"7EAB65B8",
x"7EF1659B",
x"7F4165C2",
x"7F91662A",
x"7FD966C2",
x"8010677F",
x"8032684C",
x"803B6916",
x"802F69CE",
x"80146A63",
x"7FF36ACE",
x"7FD96B0A",
x"7FD66B19",
x"7FF66B00",
x"80426AC8",
x"80C26A7D",
x"81766A30",
x"825969E9",
x"836269B8",
x"848169A6",
x"85AA69B5",
x"86CB69ED",
x"87DB6A4E",
x"88CC6AD1",
x"899B6B70",
x"8A426C26",
x"8AC26CE6",
x"8B1B6DA6",
x"8B506E57",
x"8B666EEF",
x"8B5D6F65",
x"8B3C6FAD",
x"8B076FC4",
x"8AC46FA7",
x"8A776F59",
x"8A2B6EE1",
x"89E66E4A",
x"89AB6D9E",
x"897E6CF0",
x"895F6C4E",
x"89486BC5",
x"89326B61",
x"89146B28",
x"88E46B1C",
x"889B6B37",
x"88316B72",
x"87A76BC4",
x"87036C1D",
x"864C6C73",
x"85916CB8",
x"84E06CE8",
x"84446CFA",
x"83C86CF3",
x"836F6CD4",
x"833B6CA1",
x"83246C63",
x"83236C21",
x"83286BDE",
x"832B6B9D",
x"83216B5E",
x"83016B20",
x"82CB6AE1",
x"827E6A9A",
x"82216A4B",
x"81B969F2",
x"814E698E",
x"80E26921",
x"807A68AE",
x"80146837",
x"7FAC67BC",
x"7F3C6742",
x"7EBA66C8",
x"7E1A6649",
x"7D5565C8",
x"7C62653E",
x"7B3B64AA",
x"79E0640D",
x"78556369",
x"76A062C1",
x"74D2621B",
x"72FA6181",
x"713460FC",
x"6F996093",
x"6E48604F",
x"6D606033",
x"6CFF6046",
x"6D3E6087",
x"6E3160F2",
x"6FDE6183",
x"72446237",
x"75516307",
x"78E763F2",
x"7CE264F2",
x"81106607",
x"853F6732",
x"893C6873",
x"8CDC69C9",
x"90016B35",
x"92976CB4",
x"949C6E41",
x"961F6FD4",
x"97367161",
x"980472DE",
x"98A9743D",
x"99487572",
x"99F77677",
x"9AC37744",
x"9BAE77DA",
x"9CAB783D",
x"9DA77874",
x"9E85788C",
x"9F32788F",
x"9F98788C",
x"9FAC788B",
x"9F6D7890",
x"9EE9789F",
x"9E2F78B3",
x"9D5A78C8",
x"9C8178D3",
x"9BB878CB",
x"9B0B78A9",
x"9A807862",
x"9A1177F7",
x"99B27762",
x"995976AC",
x"98F675D8",
x"988474F1",
x"98037400",
x"97787312",
x"96F6722F",
x"968B7165",
x"964D70BD",
x"9645703D",
x"967A6FEE",
x"96E66FD1",
x"97786FE8",
x"981B702D",
x"98B6709C",
x"992F7129",
x"997371C7",
x"9979726C",
x"99437309",
x"98DF7395",
x"98627405",
x"97E6745A",
x"97877493",
x"975C74BA",
x"977674D8",
x"97DC74FB",
x"988D7531",
x"99807583",
x"9AA875FC",
x"9BF37699",
x"9D4D7758",
x"9EA7782F",
x"9FEC7908",
x"A10B79D4",
x"A1F77A7B",
x"A29B7AEA",
x"A2E97B12",
x"A2D37AEB",
x"A24F7A72",
x"A15779AF",
x"9FF378AC",
x"9E2E777C",
x"9C1F7636",
x"99E774EF",
x"97AC73BE",
x"959172B6",
x"93B571E1",
x"92327148",
x"911370EE",
x"905570CA",
x"8FE670D4",
x"8FB270FF",
x"8F98713A",
x"8F7D7175",
x"8F4671A3",
x"8EEA71B9",
x"8E6571B0",
x"8DBF7188",
x"8D107143",
x"8C6F70EE",
x"8BF47093",
x"8BB67044",
x"8BBF700C",
x"8C0D6FF6",
x"8C917009",
x"8D357045",
x"8DD670A3",
x"8E537113",
x"8E8E7188",
x"8E6F71E9",
x"8DEA7229",
x"8D067237",
x"8BCF720A",
x"8A6071A3",
x"88D97103",
x"875B7037",
x"85FC6F4B",
x"84CE6E4D",
x"83D26D42",
x"82FC6C35",
x"822F6B23",
x"814B6A04",
x"802568CF",
x"7E9B6776",
x"7C8E65F2",
x"79F26439",
x"76C46250",
x"731B6042",
x"6F1D5E1E",
x"6AFC5BFE",
x"66F259FD",
x"633B5836",
x"601056C0",
x"5DA155B0",
x"5C0D550E",
x"5B6454DA",
x"5BA65511",
x"5CC455A3",
x"5EA05681",
x"61195795",
x"640358CD",
x"67375A18",
x"6A8C5B6B",
x"6DE25CBB",
x"711A5E03",
x"74235F42",
x"76EB6077",
x"796961A5",
x"7B9B62CE",
x"7D8363F3",
x"7F256517",
x"808A663A",
x"81BB675C",
x"82C56879",
x"83B26991",
x"84906A9E",
x"85656B9D",
x"86346C87",
x"87006D58",
x"87C26E08",
x"88726E92",
x"89016EF2",
x"89636F21",
x"898A6F20",
x"896D6EEB",
x"89086E83",
x"88626DEE",
x"87846D2E",
x"86806C51",
x"856D6B5C",
x"84636A5F",
x"83776965",
x"82BB687F",
x"823567B7",
x"81E6671A",
x"81C666B1",
x"81C96681",
x"81DF668D",
x"81F766CE",
x"820A673C",
x"821167CE",
x"82106872",
x"82136919",
x"822469B5",
x"82536A3B",
x"82AA6A9E",
x"832D6ADC",
x"83D56AF3",
x"84976AEB",
x"855D6AC9",
x"86106A9D",
x"86986A70",
x"86E26A4F",
x"86E36A41",
x"86A06A4B",
x"86246A72",
x"85866AB2",
x"84E66B09",
x"84656B75",
x"841D6BED",
x"84276C70",
x"848B6CFD",
x"85496D8F",
x"86506E23",
x"87886EB7",
x"88D26F47",
x"8A096FCA",
x"8B0A7039",
x"8BBF7085",
x"8C1570A7",
x"8C077094",
x"8B9B7047",
x"8ADF6FBD",
x"89EA6EFE",
x"88D66E12",
x"87BE6D0A",
x"86B56BF9",
x"85CF6AF2",
x"85136A07",
x"84836947",
x"841A68B8",
x"83CE685C",
x"83956830",
x"83626828",
x"832E683C",
x"82F3685F",
x"82B16884",
x"826D68A6",
x"822E68BC",
x"81FD68CB",
x"81E368D2",
x"81E268D5",
x"81FC68DB",
x"822B68E6",
x"826968F6",
x"82AB690A",
x"82E4691D",
x"83096928",
x"83136927",
x"82FD6910",
x"82CB68E2",
x"8284689B",
x"82316841",
x"81E067D6",
x"819B6762",
x"816966EC",
x"8149667C",
x"81386611",
x"812165AE",
x"80F0654E",
x"808A64E9",
x"7FD16476",
x"7EAC63EF",
x"7D0D634B",
x"7AEF628A",
x"785961AE",
x"756660C1",
x"723D5FCC",
x"6F095EE0",
x"6C025E0D",
x"69585D60",
x"67375CE4",
x"65BD5CA1",
x"64F95C97",
x"64E85CC2",
x"65765D18",
x"66865D8E",
x"67EF5E17",
x"69895EA4",
x"6B2B5F2B",
x"6CBB5FA4",
x"6E246007",
x"6F5B6058",
x"70656095",
x"714B60C9",
x"721D60F9",
x"72E9612F",
x"73C16177",
x"74AE61D9",
x"75B8625C",
x"76DF6303",
x"782063CC",
x"797664B4",
x"7AD965B1",
x"7C4266B4",
x"7DAA67B0",
x"7F0B6893",
x"80666951",
x"81B769E1",
x"83006A3B",
x"843F6A65",
x"85766A65",
x"86A56A47",
x"87CB6A1D",
x"88E369F7",
x"89EC69E8",
x"8ADC69F6",
x"8BAE6A28",
x"8C5C6A7F",
x"8CDF6AF0",
x"8D356B70",
x"8D5F6BF5",
x"8D5F6C6D",
x"8D416CD4",
x"8D126D21",
x"8CE56D59",
x"8CC96D82",
x"8CD36DA4",
x"8D0E6DCA",
x"8D846DFD",
x"8E356E45",
x"8F1B6EA0",
x"90296F0C",
x"91506F7F",
x"927A6FF0",
x"93987054",
x"949870A0",
x"957370D4",
x"962470EE",
x"96AC70F4",
x"971170EC",
x"975970E2",
x"978A70DF",
x"97A870E8",
x"97B670FF",
x"97B37123",
x"979E7151",
x"97747180",
x"973871AD",
x"96F071D5",
x"96A771F9",
x"9669721A",
x"964B7243",
x"96597276",
x"969F72C0",
x"97227323",
x"97DF73A0",
x"98C57433",
x"99C274D1",
x"9AB9756E",
x"9B9175FC",
x"9C32766E",
x"9C8A76B7",
x"9C9176D1",
x"9C4876B7",
x"9BB9766C",
x"9AF475F2",
x"9A0D7554",
x"99147499",
x"981773CD",
x"971D72F6",
x"96297220",
x"95387154",
x"94457096",
x"934B6FF0",
x"92496F69",
x"91456F05",
x"90496EC8",
x"8F666EB5",
x"8EAF6ECE",
x"8E396F12",
x"8E126F78",
x"8E436FFC",
x"8ECB7094",
x"8F9B7135",
x"909F71D7",
x"91BB726B",
x"92C972E8",
x"93AC7345",
x"9449737C",
x"948D7389",
x"9473736B",
x"94017323",
x"934672B6",
x"925C722B",
x"9158718D",
x"905570E4",
x"8F5D7035",
x"8E776F8A",
x"8D986EDE",
x"8CA86E2B",
x"8B876D68",
x"8A0D6C80",
x"88176B62",
x"858A69FD",
x"82596845",
x"7E8B6637",
x"7A3F63DC",
x"75A8614B",
x"71075EA8",
x"6CAA5C1F",
x"68DF59E3",
x"65EB5824",
x"6406570B",
x"634C56B3",
x"63C75729",
x"655E5861",
x"67E95A3F",
x"6B2E5C9B",
x"6EE95F3C",
x"72D561EF",
x"76B7647A",
x"7A5966B4",
x"7D9A6880",
x"806669CE",
x"82B86AA1",
x"84956B09",
x"860B6B1C",
x"872B6AFC",
x"88066AC5",
x"88AA6A97",
x"89256A86",
x"89806A9D",
x"89C36AE5",
x"89F36B58",
x"8A146BEC",
x"8A2C6C93",
x"8A416D3F",
x"8A536DDF",
x"8A676E66",
x"8A7D6ECD",
x"8A916F0D",
x"8A9D6F27",
x"8A9A6F1E",
x"8A7E6EFC",
x"8A456EC8",
x"89E46E8C",
x"895D6E4E",
x"88B26E16",
x"87E76DE5",
x"870A6DBD",
x"86286D99",
x"854F6D75",
x"84906D4D",
x"83F66D1D",
x"838A6CE2",
x"83506C9D",
x"83486C4F",
x"836D6C02",
x"83B86BBA",
x"84206B82",
x"849B6B63",
x"85246B65",
x"85B66B90",
x"86526BE5",
x"86F96C68",
x"87AF6D14",
x"887E6DE8",
x"89696ED7",
x"8A716FD9",
x"8B9A70E4",
x"8CDC71E8",
x"8E2F72DA",
x"8F8873AF",
x"90DA745A",
x"921574D2",
x"932A7517",
x"940D7525",
x"94B874FE",
x"952574A9",
x"9556742F",
x"954F739C",
x"951772FE",
x"94B97262",
x"944071D5",
x"93B97165",
x"9331711A",
x"92B270F9",
x"92457106",
x"91F47140",
x"91C671A1",
x"91BE7227",
x"91DC72C5",
x"921B7372",
x"92747425",
x"92D974CE",
x"933C7567",
x"938A75E2",
x"93B2763C",
x"93A5766A",
x"9357766E",
x"92C67644",
x"91F675F4",
x"90F3757F",
x"8FD074F2",
x"8EA77454",
x"8D9173B0",
x"8CA77312",
x"8BFD7282",
x"8B9F7203",
x"8B90719A",
x"8BC67145",
x"8C3570FF",
x"8CC370C1",
x"8D567082",
x"8DD3703B",
x"8E256FE6",
x"8E3C6F82",
x"8E126F0F",
x"8DB16E94",
x"8D256E1C",
x"8C8D6DB3",
x"8C076D68",
x"8BB86D48",
x"8BBE6D5C",
x"8C2F6DA9",
x"8D176E29",
x"8E6F6ED2",
x"901A6F92",
x"91ED704E",
x"93AC70E9",
x"95127148",
x"95D7714B",
x"95BE70DC",
x"94946FEF",
x"92456E80",
x"8ED66C9A",
x"8A6D6A54",
x"854F67CE",
x"7FD56531",
x"7A6562AD",
x"7569606C",
x"713E5E98",
x"6E305D53",
x"6C685CAF",
x"6BF35CB3",
x"6CC15D59",
x"6EA05E8B",
x"7152602E",
x"7490621F",
x"78136439",
x"7B9E665B",
x"7F066863",
x"82316A41",
x"85146BE6",
x"87B86D51",
x"8A296E85",
x"8C7B6F92",
x"8EBF7085",
x"91007170",
x"93437265",
x"958B736E",
x"97D27492",
x"9A1575D2",
x"9C52772F",
x"9E85789D",
x"A0B47A13",
x"A2E07B82",
x"A50E7CDE",
x"A7407E1B",
x"A96E7F28",
x"AB8F8002",
x"AD8B80A2",
x"AF4A8102",
x"B0B28126",
x"B1A5810F",
x"B20C80C3",
x"B1DE804C",
x"B11B7FB3",
x"AFCF7F05",
x"AE187E50",
x"AC1B7D9F",
x"AA017CFC",
x"A7F47C71",
x"A61B7C04",
x"A4977BB6",
x"A3777B85",
x"A2BF7B6E",
x"A2697B6A",
x"A2617B71",
x"A28E7B7B",
x"A2D67B84",
x"A31E7B88",
x"A3537B85",
x"A36A7B7E",
x"A35D7B75",
x"A3337B6E",
x"A2F87B6D",
x"A2B67B71",
x"A27E7B79",
x"A2577B84",
x"A24A7B88",
x"A2557B82",
x"A2707B6B",
x"A2927B40",
x"A2AE7B01",
x"A2B67AAD",
x"A2A47A50",
x"A27079EF",
x"A21F7998",
x"A1B67953",
x"A1407928",
x"A0C8791B",
x"A059792C",
x"9FFA7956",
x"9FAC798C",
x"9F6A79C3",
x"9F2979E8",
x"9EDC79F1",
x"9E7079CE",
x"9DD57979",
x"9CFE78EF",
x"9BE47836",
x"9A877752",
x"98ED7654",
x"9727754A",
x"95467441",
x"9366734A",
x"919E726E",
x"900471B5",
x"8EAF7126",
x"8DAB70BE",
x"8D03707A",
x"8CB57057",
x"8CBC704E",
x"8D0D705B",
x"8D987078",
x"8E4870A1",
x"8F0870DA",
x"8FC9711C",
x"907D716E",
x"911A71CF",
x"91A17243",
x"921872CA",
x"92887365",
x"93007413",
x"938B74D4",
x"943475A0",
x"94FD7674",
x"95E47747",
x"96E37810",
x"97EA78CA",
x"98EA796D",
x"99D679F1",
x"9A9F7A57",
x"9B437AA0",
x"9BC27ACE",
x"9C1B7AE5",
x"9C557AE7",
x"9C6C7AD6",
x"9C5A7AAD",
x"9C107A64",
x"9B7079EF",
x"9A5A7940",
x"98AE7844",
x"964F76EF",
x"932C753B",
x"8F4F7329",
x"8AD570C5",
x"85F36E2B",
x"80F66B7D",
x"7C3768E6",
x"78136694",
x"74DB64B1",
x"72D16360",
x"721862B8",
x"72B762C1",
x"748E6370",
x"776964AD",
x"7AF96655",
x"7EE7683E",
x"82E06A3B",
x"869D6C26",
x"89E36DDE",
x"8C956F4F",
x"8EAE7075",
x"903B7151",
x"915971F2",
x"9232726F",
x"92F172DC",
x"93BC7351",
x"94B473DE",
x"95E77490",
x"975F756B",
x"9915766C",
x"9AF9778F",
x"9CF778C6",
x"9EF87A08",
x"A0E67B49",
x"A2B17C7C",
x"A44A7D9E",
x"A5B27EA6",
x"A6E77F8F",
x"A7F3805A",
x"A8E18107",
x"A9C08194",
x"AA9E8200",
x"AB87824F",
x"AC828282",
x"AD9782A2",
x"AEC782B5",
x"B01282C5",
x"B17182DE",
x"B2E1830F",
x"B45C835E",
x"B5DA83D6",
x"B7538476",
x"B8C3853C",
x"BA22861F",
x"BB688714",
x"BC92880D",
x"BD9B88F9",
x"BE7F89CD",
x"BF3F8A81",
x"BFDA8B15",
x"C0548B8D",
x"C0AD8BED",
x"C0EA8C3F",
x"C1088C8D",
x"C1078CD8",
x"C0E08D20",
x"C08C8D5B",
x"C0048D7D",
x"BF408D76",
x"BE3D8D35",
x"BD018CB4",
x"BB958BED",
x"BA0F8AE9",
x"B88889B6",
x"B7228874",
x"B5FE873C",
x"B53A8632",
x"B4EE856E",
x"B5238505",
x"B5DB8500",
x"B7088559",
x"B88C8604",
x"BA4786EC",
x"BC1287F3",
x"BDC98901",
x"BF4A8A03",
x"C0848AE9",
x"C16B8BAE",
x"C1FF8C55",
x"C24E8CE3",
x"C2658D63",
x"C2548DDC",
x"C2298E4F",
x"C1E88EB8",
x"C18F8F0A",
x"C10E8F32",
x"C0538F1A",
x"BF468EAA",
x"BDD18DD5",
x"BBE78C91",
x"B9828AE6",
x"B6B088E4",
x"B38C86AC",
x"B03C8466",
x"ACF5823D",
x"A9E9805D",
x"A74D7EED",
x"A54A7E02",
x"A3FB7DA8",
x"A3697DD7",
x"A3827E7A",
x"A42C7F68",
x"A535807A",
x"A667817E",
x"A78A824A",
x"A86682BC",
x"A8D682BD",
x"A8C2824C",
x"A81F8170",
x"A6FB8040",
x"A56E7EDD",
x"A39A7D65",
x"A19F7BFB",
x"9F9E7AB3",
x"9DAE7999",
x"9BD378AD",
x"9A0877E0",
x"98357715",
x"9638762D",
x"93EC7503",
x"912B737E",
x"8DE07185",
x"8A046F14",
x"85A56C3B",
x"80EC6914",
x"7C1465CE",
x"776C629E",
x"73455FBE",
x"6FF05D69",
x"6DB35BCB",
x"6CB55B04",
x"6D0E5B22",
x"6EB05C1E",
x"71735DDF",
x"751E603E",
x"79696309",
x"7E09660E",
x"82BB6920",
x"874B6C16",
x"8B976ED8",
x"8F917158",
x"933B7395",
x"969F7599",
x"99D27774",
x"9CE47934",
x"9FE17AE8",
x"A2CF7C98",
x"A5A37E43",
x"A8577FE6",
x"AAD98177",
x"AD1582E7",
x"AF058429",
x"B09E8531",
x"B1DE85F7",
x"B2C9867B",
x"B36686C0",
x"B3BA86D2",
x"B3CD86BB",
x"B39F8688",
x"B3328646",
x"B28285FD",
x"B18C85B1",
x"B0518560",
x"AED48505",
x"AD1C8498",
x"AB3C840C",
x"A943835C",
x"A749827D",
x"A5648172",
x"A3AB8043",
x"A2307EFC",
x"A1017DB0",
x"A0247C78",
x"9F987B6B",
x"9F5A7A9D",
x"9F637A1D",
x"9FA279EF",
x"A00E7A11",
x"A0977A72",
x"A12F7B01",
x"A1C97BA2",
x"A25A7C3C",
x"A2D57CB7",
x"A32F7D02",
x"A3617D12",
x"A3667CE5",
x"A3397C82",
x"A2D97BF2",
x"A24C7B47",
x"A1987A8F",
x"A0CD79D7",
x"9FFD792A",
x"9F3B7890",
x"9E9D780C",
x"9E39779F",
x"9E247748",
x"9E69770B",
x"9F1176E5",
x"A01576DA",
x"A16D76EC",
x"A301771D",
x"A4B5776C",
x"A66A77DA",
x"A7FE7860",
x"A95678F5",
x"AA597990",
x"AAFB7A28",
x"AB387AB0",
x"AB177B20",
x"AAA87B72",
x"AA007BA8",
x"A9387BC0",
x"A8697BC6",
x"A7A97BC1",
x"A70A7BBC",
x"A6947BC0",
x"A64F7BD6",
x"A63B7BFE",
x"A6537C37",
x"A6917C7E",
x"A6ED7CC6",
x"A75C7D06",
x"A7D47D32",
x"A84F7D41",
x"A8C07D2F",
x"A9227CFB",
x"A96B7CA8",
x"A9957C41",
x"A99E7BD1",
x"A9827B68",
x"A9437B0F",
x"A8E47AD0",
x"A86A7AAC",
x"A7DA7AA3",
x"A73A7AAD",
x"A68F7ABE",
x"A5DC7ACB",
x"A51C7AC7",
x"A4507AA8",
x"A3717A6A",
x"A27D7A0C",
x"A1697995",
x"A0317909",
x"9ECF7874",
x"9D3D77D7",
x"9B737734",
x"99677686",
x"970E75C3",
x"945C74D7",
x"914073AD",
x"8DB47234",
x"89B2705B",
x"85416E1C",
x"80706B79",
x"7B636887",
x"76456562",
x"71516232",
x"6CC45F25",
x"68DE5C6C",
x"65D75A30",
x"63D9589B",
x"62FD57BF",
x"634757A5",
x"649E5845",
x"66DC5984",
x"69C55B40",
x"6D175D4C",
x"70905F78",
x"73EF619A",
x"77016386",
x"79A26524",
x"7BC46663",
x"7D5F673F",
x"7E8367C2",
x"7F4667FC",
x"7FC56804",
x"801B67F6",
x"806267E8",
x"80AA67ED",
x"81016814",
x"816A6863",
x"81E668D9",
x"826D6970",
x"82FC6A1E",
x"838A6AD8",
x"84176B90",
x"84A16C3D",
x"85286CD7",
x"85AE6D5B",
x"86356DC5",
x"86C16E19",
x"874C6E58",
x"87D66E86",
x"88566EA7",
x"88C56EBF",
x"891B6ED2",
x"89506EDF",
x"89606EE9",
x"89486EEF",
x"89086EF2",
x"88A86EEC",
x"882D6EE1",
x"87A06ECA",
x"870D6EA6",
x"867D6E76",
x"85F76E38",
x"85836DEE",
x"85216D97",
x"84D56D3D",
x"849D6CE1",
x"84766C8A",
x"845A6C3F",
x"84456C04",
x"84316BDC",
x"84186BC8",
x"83F66BC8",
x"83C86BD7",
x"838E6BEF",
x"834E6C0A",
x"830B6C23",
x"82D66C38",
x"82B86C45",
x"82BF6C4F",
x"82FC6C59",
x"83736C69",
x"842C6C86",
x"85286CB4",
x"865C6CF9",
x"87BF6D51",
x"893E6DBB",
x"8AC86E31",
x"8C4B6EA9",
x"8DB66F1A",
x"8F036F7C",
x"90286FC8",
x"91256FFC",
x"91FE7019",
x"92B47021",
x"934B7019",
x"93C27008",
x"94176FF2",
x"94406FDB",
x"94386FC5",
x"93F16FB4",
x"936A6FA3",
x"929E6F94",
x"91976F89",
x"90626F82",
x"8F156F83",
x"8DCC6F92",
x"8CA26FB5",
x"8BB46FF2",
x"8B117048",
x"8AC570B9",
x"8ACE713A",
x"8B1B71C3",
x"8B977245",
x"8C2572B1",
x"8CA872F8",
x"8D04730C",
x"8D2772E8",
x"8D077289",
x"8CA771F5",
x"8C147134",
x"8B607055",
x"8AA26F66",
x"89F06E78",
x"89596D93",
x"88E96CC1",
x"88A16C07",
x"887D6B65",
x"88706AD8",
x"886A6A5C",
x"885C69E9",
x"8832697A",
x"87E06909",
x"8758688E",
x"86906807",
x"857F676F",
x"842166C2",
x"827365FD",
x"8072651E",
x"7E22642A",
x"7B8E6323",
x"78C7620E",
x"75E560F9",
x"73065FEE",
x"704F5EFE",
x"6DE95E35",
x"6BF95D9E",
x"6A9A5D45",
x"69E35D2E",
x"69DE5D59",
x"6A825DC2",
x"6BC15E63",
x"6D7F5F33",
x"6F9B6029",
x"71F7613B",
x"7472625F",
x"76F26390",
x"796564C6",
x"7BC265FD",
x"7E066732",
x"802E685F",
x"823C6980",
x"84346A90",
x"86136B8A",
x"87D96C6D",
x"89806D35",
x"8B036DE5",
x"8C5D6E7F",
x"8D8E6F09",
x"8E926F88",
x"8F6D7002",
x"90247080",
x"90B87105",
x"91327195",
x"9194722D",
x"91E072CD",
x"9214736F",
x"9231740D",
x"923274A1",
x"92177523",
x"91E0758D",
x"919175DB",
x"91317609",
x"90CB7615",
x"906A7602",
x"901D75D2",
x"8FEE758C",
x"8FED7539",
x"901F74E2",
x"908D7495",
x"9135745E",
x"9218744B",
x"93347468",
x"948074C0",
x"95FA7555",
x"979B762D",
x"995F7746",
x"9B3C7898",
x"9D2C7A18",
x"9F247BB7",
x"A1157D65",
x"A2F37F0B",
x"A4A98098",
x"A62B81F7",
x"A7668317",
x"A85083E8",
x"A8E78467",
x"A92F848F",
x"A9338467",
x"A90883FA",
x"A8CC835A",
x"A89C82A2",
x"A89E81EE",
x"A8F1815B",
x"A9B58107",
x"AAFE810A",
x"ACDA8177",
x"AF4D8259",
x"B25383B3",
x"B5DE857E",
x"B9D487AC",
x"BE168A27",
x"C2818CD2",
x"C6E88F8E",
x"CB23923F",
x"CF0994C5",
x"D2749702",
x"D54698DF",
x"D7679A4A",
x"D8C89B33",
x"D9689B93",
x"D94A9B69",
x"D87E9ABA",
x"D716998F",
x"D52C97F9",
x"D2DA960F",
x"D03993E9",
x"CD6791A8",
x"CA7C8F6A",
x"C7958D50",
x"C4CA8B76",
x"C23589F4",
x"BFEE88DC",
x"BE0B8835",
x"BC998800",
x"BBA2882F",
x"BB2288AF",
x"BB0B8963",
x"BB428A2B",
x"BBA58AE6",
x"BC0B8B74",
x"BC478BBC",
x"BC388BAF",
x"BBBC8B48",
x"BAC98A88",
x"B9608983",
x"B791884C",
x"B57886FB",
x"B33C85AE",
x"B0FE8477",
x"AEDE8366",
x"ACF1827E",
x"AB3281B7",
x"A9948102",
x"A7F48042",
x"A6257F56",
x"A3F47E20",
x"A1307C82",
x"9DB57A6A",
x"996C77D2",
x"945774C3",
x"8E917152",
x"884C6DA6",
x"81CF69E6",
x"7B696649",
x"757062FA",
x"70376025",
x"6C005DE7",
x"68FB5C50",
x"67415B67",
x"66D15B21",
x"67945B6B",
x"69615C2E",
x"6BFF5D4B",
x"6F355EAB",
x"72C56035",
x"767C61DA",
x"7A2B638B",
x"7DB46542",
x"80FE66F7",
x"840368A6",
x"86BE6A47",
x"89326BD4",
x"8B666D45",
x"8D606E96",
x"8F2B6FC0",
x"90CF70C1",
x"925671A0",
x"93CB7264",
x"9538731A",
x"96A773D2",
x"9821749C",
x"99AB7581",
x"9B487689",
x"9CF377B2",
x"9EA278F2",
x"A0487A39",
x"A1D07B6F",
x"A3287C7C",
x"A43D7D49",
x"A4FE7DC0",
x"A5637DD6",
x"A5667D89",
x"A50B7CE1",
x"A45A7BEF",
x"A3647ACB",
x"A2387992",
x"A0EA785E",
x"9F8B774A",
x"9E2C766B",
x"9CDC75CB",
x"9BA57572",
x"9A91755A",
x"99A57578",
x"98E775C1",
x"98597623",
x"97FA768F",
x"97C976F7",
x"97C0774D",
x"97D87788",
x"980377A3",
x"9833779C",
x"985A776E",
x"9869771D",
x"985076AD",
x"980A761F",
x"9790757C",
x"96E774CB",
x"96187416",
x"952F7366",
x"943F72C5",
x"9359723B",
x"928E71CF",
x"91ED7183",
x"917E715B",
x"91487151",
x"91467165",
x"91777190",
x"91D571D1",
x"92567223",
x"92F37288",
x"93A772FE",
x"946D738C",
x"95437436",
x"962C74FC",
x"972775E0",
x"983576DD",
x"995677EB",
x"9A8878FB",
x"9BC879FB",
x"9D0D7AD8",
x"9E4A7B82",
x"9F767BE5",
x"A07D7BF9",
x"A1527BBD",
x"A1E97B39",
x"A2387A79",
x"A23D7998",
x"A20178B2",
x"A18F77E4",
x"A103774B",
x"A0777703",
x"A00F7718",
x"9FED7790",
x"A02B786A",
x"A0D97993",
x"A1FD7AF8",
x"A38A7C7C",
x"A5677E02",
x"A7707F6D",
x"A97580A6",
x"AB4F81A1",
x"ACD28250",
x"ADE082B8",
x"AE6E82DD",
x"AE7D82CC",
x"AE198294",
x"AD618243",
x"AC7781E8",
x"AB76818C",
x"AA788133",
x"A98E80DB",
x"A8B6807E",
x"A7E1800E",
x"A6F47F7E",
x"A5CA7EBC",
x"A43F7DB7",
x"A22B7C61",
x"9F777AB2",
x"9C1578A3",
x"9808763D",
x"9369738B",
x"8E5A70A0",
x"89136D9A",
x"83CC6A9A",
x"7EC667C2",
x"7A3F6537",
x"766C6313",
x"7375616F",
x"71726059",
x"706F5FD3",
x"70625FD8",
x"71386056",
x"72CF6137",
x"74FF625F",
x"779B63B4",
x"7A7C6520",
x"7D79668B",
x"807367EF",
x"83506941",
x"86046A84",
x"88846BBF",
x"8ACE6CF9",
x"8CE06E3B",
x"8EC16F8C",
x"907370EF",
x"91F9725E",
x"935373D2",
x"9481753A",
x"957D7685",
x"9646779D",
x"96D77872",
x"972F78F8",
x"97507928",
x"97427908",
x"971078A5",
x"96CC7815",
x"96887778",
x"965D76EB",
x"965D768C",
x"969A7672",
x"971B76AC",
x"97E27739",
x"98E0780B",
x"9A07790E",
x"9B3C7A1F",
x"9C647B22",
x"9D667BF5",
x"9E327C85",
x"9EC27CC7",
x"9F1E7CC4",
x"9F5A7C8E",
x"9F947C44",
x"9FEE7C09",
x"A08D7C05",
x"A1887C53",
x"A2F37D08",
x"A4C97E26",
x"A6FA7FA3",
x"A96A8168",
x"ABEE8352",
x"AE5D8536",
x"B08C86F1",
x"B25D8862",
x"B3BA8973",
x"B4A18A1A",
x"B5168A5D",
x"B5358A48",
x"B51589F4",
x"B4DC897E",
x"B4A98903",
x"B49E889E",
x"B4CE886A",
x"B5508879",
x"B62988D8",
x"B75B898A",
x"B8E18A93",
x"BAAD8BE5",
x"BCAC8D74",
x"BEC18F28",
x"C0D090E7",
x"C2B49293",
x"C451940C",
x"C5899537",
x"C64695FF",
x"C67E9659",
x"C6369645",
x"C57E95D1",
x"C4729510",
x"C3389424",
x"C1F1932A",
x"C0C3923E",
x"BFC39174",
x"BEFA90D3",
x"BE5E9056",
x"BDDB8FEC",
x"BD508F79",
x"BC958EE5",
x"BB888E14",
x"BA138CFA",
x"B8328B97",
x"B5F089F9",
x"B374883B",
x"B0EE8684",
x"AE9E84FE",
x"ACC283D0",
x"AB888315",
x"AB1882DD",
x"AB788323",
x"AC9B83D4",
x"AE5384D0",
x"B06785EA",
x"B28B86F6",
x"B47387CA",
x"B5DB8845",
x"B6928854",
x"B67E87F4",
x"B59E872C",
x"B4088612",
x"B1E784C2",
x"AF71835A",
x"ACDD81F6",
x"AA5480A9",
x"A7F57F7C",
x"A5C37E70",
x"A3AC7D6D",
x"A1877C5A",
x"9F197B13",
x"9C287977",
x"98797760",
x"93E774BA",
x"8E67717F",
x"880A6DB8",
x"81036986",
x"79A26518",
x"724F60AD",
x"6B765C86",
x"658258E4",
x"60CC5602",
x"5D975405",
x"5C0252FF",
x"5C0652ED",
x"5D7F53B3",
x"602D552B",
x"63C05721",
x"67DE5960",
x"6C345BB9",
x"707C5E06",
x"747D602B",
x"7817621E",
x"7B3863DA",
x"7DE26569",
x"801B66CE",
x"81F36810",
x"83766932",
x"84AF6A32",
x"85A46B09",
x"86556BB0",
x"86C36C1E",
x"86F06C55",
x"86E06C55",
x"869D6C2A",
x"86356BE2",
x"85BC6B8F",
x"85486B44",
x"84EA6B0D",
x"84B46AF5",
x"84AC6AFD",
x"84D66B21",
x"852A6B58",
x"859B6B93",
x"86186BC4",
x"86936BE3",
x"86FC6BE8",
x"87496BD2",
x"877A6BA6",
x"87916B6B",
x"87966B2B",
x"87946AF0",
x"87986AC4",
x"87AB6AAA",
x"87D26AA4",
x"880B6AB1",
x"884F6ACB",
x"88936AEF",
x"88C66B16",
x"88D86B3B",
x"88BC6B5C",
x"88696B76",
x"87DB6B8D",
x"87186BA0",
x"862C6BB2",
x"852B6BC7",
x"84276BDC",
x"83376BF5",
x"826D6C0D",
x"81DB6C26",
x"81846C38",
x"816A6C41",
x"81846C3E",
x"81C66C2B",
x"821B6C07",
x"82736BD2",
x"82BC6B8D",
x"82E96B3B",
x"82EF6AE1",
x"82CF6A80",
x"82896A20",
x"822569C1",
x"81AE6965",
x"812D690D",
x"80AD68B7",
x"80346860",
x"7FC86807",
x"7F6967AA",
x"7F17674B",
x"7ECE66EB",
x"7E876691",
x"7E3E6646",
x"7DEF6617",
x"7D95660B",
x"7D346630",
x"7CC96686",
x"7C5E6711",
x"7BF767CC",
x"7BA068AB",
x"7B5F699E",
x"7B3E6A91",
x"7B426B6F",
x"7B6F6C24",
x"7BC26C9E",
x"7C386CD8",
x"7CC96CCE",
x"7D6A6C86",
x"7E116C12",
x"7EB46B82",
x"7F4E6AED",
x"7FDC6A6C",
x"80606A13",
x"80E069EC",
x"81656A02",
x"81F26A4F",
x"82916ACF",
x"83426B72",
x"84066C24",
x"84D56CD4",
x"85A26D6F",
x"86606DE8",
x"87016E33",
x"87746E4D",
x"87AC6E33",
x"879E6DE6",
x"87436D6C",
x"86976CC7",
x"85936BF6",
x"84376AFD",
x"828069D9",
x"80706889",
x"7E09670A",
x"7B53655F",
x"785D6390",
x"753B61A5",
x"720C5FB1",
x"6EF05DC8",
x"6C135C02",
x"69995A7A",
x"67A95943",
x"665C5870",
x"65C5580C",
x"65E5581C",
x"66AE589B",
x"6809597D",
x"69CF5AAE",
x"6BDB5C1B",
x"6E035DAC",
x"70215F4B",
x"721D60DF",
x"73E36256",
x"756C63A3",
x"76BC64BA",
x"77E26598",
x"78E9663C",
x"79E666AD",
x"7AE666F0",
x"7BF66717",
x"7D19672D",
x"7E4B6742",
x"7F816763",
x"80B1679D",
x"81C667F2",
x"82B76863",
x"837468ED",
x"83FD6986",
x"84536A20",
x"84816AB0",
x"84986B2B",
x"84AF6B89",
x"84DD6BC8",
x"85386BED",
x"85CE6C02",
x"86A86C10",
x"87C86C28",
x"891F6C58",
x"8A9D6CA8",
x"8C286D21",
x"8DA46DC4",
x"8EF66E8A",
x"90086F70",
x"90CC7066",
x"913B7164",
x"91587257",
x"912F7334",
x"90D373EF",
x"9059747F",
x"8FD874DA",
x"8F6274FB",
x"8F0774E2",
x"8ED07490",
x"8EC1740F",
x"8ED57366",
x"8F0472A9",
x"8F4271E8",
x"8F807137",
x"8FB270A7",
x"8FCC704A",
x"8FC37023",
x"8F957035",
x"8F43707C",
x"8ED070E6",
x"8E467164",
x"8DB271DF",
x"8D247245",
x"8CAA7286",
x"8C537299",
x"8C2A727E",
x"8C35723D",
x"8C7771E1",
x"8CEC717F",
x"8D8D7129",
x"8E4C70EF",
x"8F1E70DE",
x"8FF070FC",
x"90B9714B",
x"916D71C1",
x"92077255",
x"928572F8",
x"92EC739C",
x"933E7434",
x"938574BA",
x"93CC752A",
x"94157585",
x"946A75CD",
x"94C8760B",
x"952E7641",
x"95957675",
x"95F376A6",
x"963D76D2",
x"966A76F2",
x"966D76FC",
x"964176E8",
x"95E076AF",
x"954F7648",
x"949575B6",
x"93BE74FC",
x"92D67426",
x"91F37343",
x"91217262",
x"90737197",
x"8FF370F2",
x"8FA8707E",
x"8F907040",
x"8FA57039",
x"8FDD705F",
x"902770AA",
x"90707106",
x"90A47165",
x"90B571B5",
x"909571EB",
x"903F71FE",
x"8FB271EB",
x"8EF371B4",
x"8E0A7161",
x"8CFE70F9",
x"8BD97082",
x"8A9A7000",
x"893C6F75",
x"87B46ED9",
x"85EF6E23",
x"83DA6D44",
x"81636C2E",
x"7E806ADB",
x"7B346945",
x"77906773",
x"73BB6576",
x"6FEB6369",
x"6C5F6170",
x"695F5FB2",
x"672B5E52",
x"65F95D70",
x"65E65D1E",
x"66F95D62",
x"69195E2E",
x"6C145F6C",
x"6FAA60F7",
x"738C62AD",
x"776F6462",
x"7B1365FC",
x"7E4C6766",
x"8103689A",
x"833C699E",
x"850B6A80",
x"86976B57",
x"88066C33",
x"897C6D21",
x"8B106E2A",
x"8CCB6F43",
x"8EA4705E",
x"90817165",
x"92457240",
x"93C672D8",
x"94EA7325",
x"959A7321",
x"95CD72DA",
x"958D7262",
x"94F071D8",
x"9417715B",
x"93277106",
x"924370F2",
x"918D7129",
x"911871AD",
x"90F37274",
x"911B736A",
x"91877478",
x"92297583",
x"92ED7678",
x"93C07744",
x"949177DE",
x"95557841",
x"96017872",
x"96947877",
x"970E7857",
x"9771781B",
x"97C077C8",
x"98007765",
x"983176F2",
x"98567675",
x"987475F1",
x"988F756E",
x"98AB74F4",
x"98CF7492",
x"99037452",
x"994F7443",
x"99B8746E",
x"9A4374D5",
x"9AED7578",
x"9BAF764A",
x"9C7D773A",
x"9D467832",
x"9DFA7915",
x"9E8479CB",
x"9ED97A41",
x"9EEE7A6B",
x"9EC67A43",
x"9E6479D0",
x"9DDC7923",
x"9D407856",
x"9CA97782",
x"9C2E76C3",
x"9BE07633",
x"9BCB75E1",
x"9BEE75D5",
x"9C43760F",
x"9CBB7681",
x"9D3B7716",
x"9DA977B9",
x"9DED784B",
x"9DED78B4",
x"9D9B78E2",
x"9CF178C8",
x"9BF37861",
x"9AAF77B4",
x"993976D1",
x"97AE75CD",
x"962974C0",
x"94C673CA",
x"939B7300",
x"92B57279",
x"921B7241",
x"91CC725E",
x"91BE72C8",
x"91E77374",
x"9239744B",
x"92AA7539",
x"93347625",
x"93D576FC",
x"949277AF",
x"95737834",
x"9680788F",
x"97BB78C3",
x"992478DB",
x"9AAF78E4",
x"9C4B78E8",
x"9DD678EE",
x"9F3278F8",
x"A03C7901",
x"A0D67901",
x"A0EB78EB",
x"A07378B6",
x"9F767858",
x"9E0577D0",
x"9C42771F",
x"9A50764B",
x"984F7565",
x"965A7476",
x"9481738C",
x"92C072AA",
x"910771D2",
x"8F3B70F9",
x"8D397013",
x"8AE06F0C",
x"881D6DD2",
x"84E76C59",
x"814E6A9C",
x"7D7368A1",
x"798C667A",
x"75D66445",
x"729A6224",
x"7013603E",
x"6E6F5EB5",
x"6DC95DA5",
x"6E215D21",
x"6F625D29",
x"71615DB6",
x"73E85EAF",
x"76BB5FFC",
x"79A4617A",
x"7C7A6310",
x"7F2264A8",
x"81966635",
x"83D967B5",
x"86016928",
x"88286A9C",
x"8A636C19",
x"8CC66DA9",
x"8F596F4E",
x"92157108",
x"94EF72CA",
x"97CF7488",
x"9A9B762F",
x"9D3B77AC",
x"9F9978F2",
x"A1A979F9",
x"A3667AC3",
x"A4D27B57",
x"A5F77BC7",
x"A6E47C25",
x"A7AE7C86",
x"A8617CFF",
x"A9147D9C",
x"A9D37E63",
x"AAA87F51",
x"AB9E8064",
x"ACB9818A",
x"ADF882B3",
x"AF5E83CF",
x"B0E184CF",
x"B27885A5",
x"B417864F",
x"B5AC86C8",
x"B7288714",
x"B87A8739",
x"B995873F",
x"BA71872B",
x"BB0C8705",
x"BB6B86D3",
x"BB998699",
x"BBA6865C",
x"BBA5861E",
x"BBA885E4",
x"BBC085B2",
x"BBF7858E",
x"BC4D857A",
x"BCB98577",
x"BD298584",
x"BD828599",
x"BDA685AF",
x"BD7485B6",
x"BCD185A1",
x"BBB0855E",
x"BA0C84E3",
x"B7F4842B",
x"B5898336",
x"B2FA8212",
x"B07E80D3",
x"AE537F94",
x"ACB57E75",
x"ABCC7D96",
x"ABB67D14",
x"AC777D02",
x"ADFA7D6B",
x"B0157E4F",
x"B28C7F9C",
x"B519813D",
x"B774830E",
x"B95D84E7",
x"BAA386A5",
x"BB298821",
x"BAE88940",
x"B9EE89F0",
x"B85B8A27",
x"B65989E7",
x"B415893C",
x"B1BD8838",
x"AF7886ED",
x"AD608574",
x"AB8583E3",
x"A9EA824A",
x"A88B80BA",
x"A7607F40",
x"A65D7DE3",
x"A5767CA3",
x"A49F7B88",
x"A3D77A93",
x"A31779C6",
x"A25D791F",
x"A1A878A2",
x"A0F77848",
x"A048780F",
x"9F9477EF",
x"9ED677DB",
x"9E0777C8",
x"9D2177A6",
x"9C1F7767",
x"9AFD76FF",
x"99BE766B",
x"986275AA",
x"96F374C3",
x"957B73C3",
x"940872BB",
x"92AA71C1",
x"916F70E4",
x"90627033",
x"8F8B6FB4",
x"8EE96F68",
x"8E746F41",
x"8E1B6F2D",
x"8DBF6F16",
x"8D3E6EDE",
x"8C706E6B",
x"8B2F6DAA",
x"89596C8D",
x"86D96B10",
x"83AD693B",
x"7FDF671D",
x"7B9364D0",
x"76FD6276",
x"7261602D",
x"6E045E15",
x"6A345C4F",
x"672E5AED",
x"65265A01",
x"64385991",
x"6468599B",
x"65A45A14",
x"67C55AF0",
x"6A935C17",
x"6DCB5D76",
x"712E5EF4",
x"747F607C",
x"778761F9",
x"7A28635D",
x"7C4B64A0",
x"7DED65B8",
x"7F1B66AA",
x"7FE96777",
x"80746827",
x"80DD68C4",
x"81416958",
x"81B769E9",
x"82526A7F",
x"831B6B1D",
x"84156BBF",
x"85366C62",
x"86746D02",
x"87BC6D92",
x"88FA6E0C",
x"8A1D6E66",
x"8B146E9D",
x"8BD56EAD",
x"8C5C6E94",
x"8CA86E58",
x"8CBF6DFF",
x"8CAB6D93",
x"8C776D20",
x"8C316CAE",
x"8BE66C4F",
x"8BA16C0C",
x"8B696BED",
x"8B466BFC",
x"8B396C3D",
x"8B446CB0",
x"8B666D52",
x"8B9A6E19",
x"8BDF6EFA",
x"8C2E6FE6",
x"8C8170CD",
x"8CD3719D",
x"8D1E7247",
x"8D5B72C1",
x"8D867306",
x"8D9A7315",
x"8D9A72F4",
x"8D8472AD",
x"8D607250",
x"8D3271EB",
x"8D00718A",
x"8CCF713D",
x"8CA47109",
x"8C8070EF",
x"8C6270EF",
x"8C4670FF",
x"8C2B7114",
x"8C0A7126",
x"8BE07126",
x"8BAE710D",
x"8B7470D7",
x"8B38707E",
x"8AFE7008",
x"8ACE6F78",
x"8AAA6ED7",
x"8A936E2E",
x"8A8A6D86",
x"8A8A6CE9",
x"8A8A6C5C",
x"8A836BE8",
x"8A6C6B8C",
x"8A3E6B4C",
x"89F76B28",
x"89986B1E",
x"89256B28",
x"88A76B42",
x"88226B65",
x"87A26B8A",
x"872C6BAB",
x"86C16BC4",
x"865F6BD2",
x"86036BD5",
x"85A46BCE",
x"853B6BC1",
x"84C26BB1",
x"84346BA6",
x"83906BA0",
x"82D66BA1",
x"820D6BA8",
x"813B6BAD",
x"80666BA8",
x"7F946B8D",
x"7EC66B54",
x"7E006AEF",
x"7D3B6A5E",
x"7C74699C",
x"7BA768B0",
x"7ACB67A1",
x"79DF667F",
x"78E56558",
x"77DF643B",
x"76D66334",
x"75D6624C",
x"74EC618A",
x"742160EC",
x"7382606D",
x"73106008",
x"72CE5FB3",
x"72B25F6A",
x"72AD5F22",
x"72A75ED6",
x"72875E81",
x"722E5E1F",
x"717D5DAC",
x"705C5D22",
x"6EB85C7D",
x"6C8C5BB6",
x"69DC5ACC",
x"66BE59BC",
x"6354588A",
x"5FCF573C",
x"5C6555E4",
x"59525494",
x"56D15363",
x"5510526A",
x"543351C4",
x"544A5182",
x"555251B0",
x"57335254",
x"59C45363",
x"5CCD54CD",
x"60135677",
x"63585840",
x"66665A07",
x"69135BAB",
x"6B445D14",
x"6CEE5E2E",
x"6E145EF0",
x"6ECE5F60",
x"6F345F8A",
x"6F665F7D",
x"6F835F53",
x"6FA45F21",
x"6FD85EF8",
x"702A5EEA",
x"70945EFA",
x"71105F27",
x"71905F6A",
x"72035FB8",
x"725B6001",
x"728D603C",
x"7294605D",
x"72726062",
x"722A604B",
x"71C8601E",
x"71595FE4",
x"70ED5FAB",
x"70905F7D",
x"704B5F63",
x"70275F66",
x"70265F87",
x"70455FC5",
x"70836018",
x"70D5607D",
x"713760E7",
x"71A06150",
x"720961B1",
x"72706200",
x"72D5623C",
x"73346264",
x"7390627A",
x"73EC627E",
x"74476277",
x"74A16269",
x"74FC6259",
x"7555624C",
x"75A86246",
x"75F56248",
x"76346252",
x"76666262",
x"76896272",
x"769B627D",
x"769E627C",
x"76946269",
x"767F623F",
x"76606200",
x"763E61AD",
x"761B6149",
x"75F960E2",
x"75DC607E",
x"75C6602B",
x"75BA5FF2",
x"75B85FD8",
x"75C15FDF",
x"75D56007",
x"75F36048",
x"761A609B",
x"764460F6",
x"76706152",
x"769D61AB",
x"76C561FD",
x"76EC624E",
x"770E62A4",
x"77306306",
x"7751637F",
x"77776414",
x"77A864C8",
x"77E66597",
x"7837667C",
x"789D6765",
x"791A6845",
x"79AE690C",
x"7A5869A7",
x"7B136A0D",
x"7BDC6A38",
x"7CAB6A2A",
x"7D7A69EB",
x"7E416987",
x"7EF96913",
x"7FA068A0",
x"80326844",
x"80B26811",
x"81256816",
x"81916859",
x"81FD68E1",
x"827269A4",
x"82F46A9A",
x"83866BB1",
x"84246CD4",
x"84C46DE9",
x"855B6ED7",
x"85D36F85",
x"86206FE1",
x"862E6FDE",
x"85F66F7C",
x"85766EC4",
x"84B16DC4",
x"83B96C99",
x"82A36B5F",
x"81816A32",
x"806C692B",
x"7F6C685B",
x"7E8467C2",
x"7DA8675B",
x"7CBE670B",
x"7BA766BA",
x"7A3D6642",
x"78606589",
x"75FD6476",
x"730D6301",
x"6FA46135",
x"6BE95F25",
x"68165CF8",
x"646F5ADC",
x"614058FE",
x"5EC55788",
x"5D31569B",
x"5CA05646",
x"5D0C5688",
x"5E5C5750",
x"605F587E",
x"62D559ED",
x"657A5B71",
x"680F5CE4",
x"6A625E27",
x"6C525F25",
x"6DD55FD6",
x"6EF06041",
x"6FB8606E",
x"704C6077",
x"70CC6070",
x"714F606C",
x"71EB607E",
x"72A460B2",
x"7378610A",
x"745B6184",
x"753B621A",
x"760962BE",
x"76B56365",
x"77346401",
x"7786648D",
x"77AB6500",
x"77AE6556",
x"779A6593",
x"777C65B8",
x"775F65C9",
x"774B65CE",
x"774865C8",
x"775865BC",
x"777C65AD",
x"77B16598",
x"77F76581",
x"784E6568",
x"78B4654C",
x"792A6534",
x"79AF6523",
x"7A48651E",
x"7AEF652D",
x"7BA46550",
x"7C62658D",
x"7D2565E5",
x"7DE36653",
x"7E9866D3",
x"7F3E6762",
x"7FD167F6",
x"804E688A",
x"80B7691B",
x"811169A8",
x"81636A2D",
x"81B46AAA",
x"82096B1E",
x"82696B8C",
x"82D66BED",
x"83526C42",
x"83D96C86",
x"84656CB8",
x"84F06CD4",
x"85766CDB",
x"85F36CD2",
x"86656CBE",
x"86D16CA7",
x"873C6C94",
x"87B56C8F",
x"88436C9A",
x"88F46CB7",
x"89CF6CE6",
x"8AD86D23",
x"8C0B6D65",
x"8D626DAA",
x"8ECB6DEB",
x"90326E26",
x"91836E5C",
x"92A46E92",
x"93816EC8",
x"940E6F06",
x"94426F4B",
x"941C6F96",
x"93A56FDE",
x"92EA701A",
x"91FB703E",
x"90EE703B",
x"8FD87009",
x"8EC66FA1",
x"8DC86F09",
x"8CE66E48",
x"8C276D73",
x"8B896C9E",
x"8B0D6BE3",
x"8AB26B59",
x"8A766B10",
x"8A596B0F",
x"8A5C6B57",
x"8A816BD9",
x"8AC96C86",
x"8B346D44",
x"8BBE6DF9",
x"8C606E8F",
x"8D116EF0",
x"8DBE6F17",
x"8E556EFE",
x"8EC16EAA",
x"8EED6E27",
x"8ECC6D85",
x"8E506CD2",
x"8D7B6C21",
x"8C556B7C",
x"8AEC6AEC",
x"895C6A79",
x"87C26A24",
x"863969EC",
x"84DA69CB",
x"83B469BA",
x"82C569AB",
x"81FE698E",
x"81436954",
x"806D68E5",
x"7F4E682E",
x"7DBB6723",
x"7B9465B7",
x"78C963EC",
x"755E61CC",
x"716C5F72",
x"6D245CFD",
x"68CA5A95",
x"64A05869",
x"60EF569E",
x"5DF55556",
x"5BDB54A3",
x"5AB6548E",
x"5A805508",
x"5B1F55F7",
x"5C675736",
x"5E1E589E",
x"600F5A04",
x"62055B43",
x"63D75C42",
x"65685CF3",
x"66AD5D52",
x"67A55D67",
x"68595D43",
x"68D85CF8",
x"692D5C9C",
x"69695C3F",
x"69945BED",
x"69B75BAF",
x"69D65B8A",
x"69F65B7B",
x"6A1D5B84",
x"6A525BA4",
x"6A9C5BD7",
x"6B035C1F",
x"6B8E5C7A",
x"6C3F5CE6",
x"6D115D62",
x"6DFD5DE6",
x"6EF25E6E",
x"6FDE5EF3",
x"70B15F6A",
x"71595FD0",
x"71D26022",
x"72186060",
x"7237608E",
x"723D60B8",
x"723E60E4",
x"72536121",
x"728D6174",
x"72F961E4",
x"7398626D",
x"7468630A",
x"755563AD",
x"764B6446",
x"773164C8",
x"77ED6523",
x"786D654E",
x"78A86548",
x"789D6513",
x"785564BB",
x"77E06452",
x"775863E9",
x"76D46394",
x"76696363",
x"762D6360",
x"7627638E",
x"765B63EC",
x"76C5646D",
x"77596504",
x"7807659B",
x"78BF6623",
x"79736689",
x"7A1466C4",
x"7A9D66CC",
x"7B0A66A4",
x"7B606656",
x"7BA465EF",
x"7BE06580",
x"7C1D6520",
x"7C6364DF",
x"7CBA64CE",
x"7D2164F3",
x"7D9A6552",
x"7E1E65E3",
x"7EA56697",
x"7F22675C",
x"7F8C681B",
x"7FD568BF",
x"7FF46934",
x"7FE7696C",
x"7FAA6961",
x"7F3F6916",
x"7EB16897",
x"7E0767F3",
x"7D526741",
x"7C9B6694",
x"7BF06600",
x"7B596594",
x"7ADC6555",
x"7A7C6545",
x"7A32655B",
x"79FF658A",
x"79D865C4",
x"79BB65F6",
x"79A46613",
x"79936611",
x"798D65EA",
x"799765A4",
x"79BA6544",
x"79FF64DA",
x"7A6A6477",
x"7AFC642A",
x"7BAD63FF",
x"7C736401",
x"7D3A6434",
x"7DF06491",
x"7E816510",
x"7EDC65A0",
x"7EF76630",
x"7ED266B0",
x"7E726710",
x"7DE36749",
x"7D386756",
x"7C816738",
x"7BCC66F7",
x"7B21669B",
x"7A7A662E",
x"79CF65B8",
x"7910653E",
x"782864BF",
x"770A6439",
x"75B163AD",
x"741E6311",
x"72686268",
x"70AE61B4",
x"6F1D6100",
x"6DE3605C",
x"6D305FD9",
x"6D275F8E",
x"6DE25F8E",
x"6F655FE9",
x"71A360A5",
x"747C61C6",
x"77C86341",
x"7B566503",
x"7EF666F6",
x"82836900",
x"85DF6B09",
x"88FC6CF6",
x"8BD96EBA",
x"8E847048",
x"911071A0",
x"938E72C5",
x"961573C4",
x"98B474AA",
x"9B707589",
x"9E4A7674",
x"A13E7778",
x"A43D78A0",
x"A73C79F7",
x"AA307B77",
x"AD0D7D1E",
x"AFC97EDD",
x"B26080A5",
x"B4CC8263",
x"B7088402",
x"B9128571",
x"BAE786A1",
x"BC87878E",
x"BDF28838",
x"BF2F88A9",
x"C04688F6",
x"C142892F",
x"C230896D",
x"C32289C3",
x"C4208A42",
x"C5368AEC",
x"C6618BBE",
x"C79C8CAE",
x"C8DE8DAA",
x"CA188E9E",
x"CB3A8F7A",
x"CC3C9031",
x"CD1890BF",
x"CDD49127",
x"CE7F9174",
x"CF2A91B8",
x"CFEF9204",
x"D0E2926A",
x"D21392F4",
x"D38B93AA",
x"D53E9483",
x"D7209578",
x"D9109676",
x"DAEE976B",
x"DC929841",
x"DDDB98E8",
x"DEB09955",
x"DF01997F",
x"DECB9966",
x"DE1A990F",
x"DD029885",
x"DB9D97D2",
x"DA0E970A",
x"D871963F",
x"D6E89589",
x"D58B94FC",
x"D46C94AA",
x"D39894A4",
x"D31094F3",
x"D2D09597",
x"D2C99684",
x"D2E297A4",
x"D30598D4",
x"D31099EC",
x"D2E49AC2",
x"D2629B30",
x"D1799B17",
x"D0199A6B",
x"CE41992D",
x"CBFC9775",
x"C9619565",
x"C689932A",
x"C39690F4",
x"C0A58EEF",
x"BDCA8D34",
x"BB188BD2",
x"B8918AC0",
x"B62E89EA",
x"B3E4892E",
x"B1A28862",
x"AF5A8764",
x"AD05861B",
x"AAA1847E",
x"A8388295",
x"A5DE807B",
x"A3AE7E59",
x"A1BF7C57",
x"A02B7AA5",
x"9F037965",
x"9E4A78AD",
x"9E017881",
x"9E1278D1",
x"9E66797F",
x"9EDD7A64",
x"9F577B4D",
x"9FB97C11",
x"9FEC7C8B",
x"9FE37CA3",
x"9F997C53",
x"9F197BA3",
x"9E6C7AAC",
x"9DA1798B",
x"9CC97862",
x"9BEE7755",
x"9B15767B",
x"9A3575DE",
x"993C7579",
x"980F753A",
x"968B74FC",
x"948A7497",
x"91E773DF",
x"8E8872AA",
x"8A5F70DB",
x"856F6E68",
x"7FD66B58",
x"79C567C8",
x"738363ED",
x"6D666006",
x"67CA5C5C",
x"63095935",
x"5F7556D0",
x"5D45555A",
x"5C9C54ED",
x"5D785582",
x"5FB75704",
x"6320593F",
x"675F5BF7",
x"6C145EE4",
x"70E161C5",
x"7569645A",
x"79656679",
x"7CA36809",
x"7F0A6906",
x"809B697D",
x"816C698E",
x"81A2695F",
x"816F6919",
x"810468E3",
x"809068DB",
x"80376911",
x"8010698A",
x"802A6A38",
x"80816B0A",
x"810D6BE2",
x"81BC6CA6",
x"827D6D3D",
x"833F6D93",
x"83F66DA4",
x"849B6D73",
x"852C6D0D",
x"85AE6C87",
x"86256BF9",
x"869A6B7D",
x"87116B24",
x"878E6AFD",
x"880D6B0C",
x"88866B49",
x"88EF6BAA",
x"893C6C1E",
x"89666C90",
x"89626CEE",
x"89326D2B",
x"88DC6D41",
x"886D6D30",
x"87F96D00",
x"87946CBF",
x"87536C80",
x"87496C54",
x"87836C4D",
x"88046C73",
x"88C86CCF",
x"89C26D5E",
x"8AE06E14",
x"8C0B6EE4",
x"8D2C6FBA",
x"8E2E7082",
x"8F017127",
x"8F9D719C",
x"8FFC71D7",
x"902171D7",
x"901771A1",
x"8FE67143",
x"8F9B70CD",
x"8F417052",
x"8EE36FE8",
x"8E876F9C",
x"8E356F79",
x"8DF16F89",
x"8DBC6FCA",
x"8D9C7035",
x"8D9470C5",
x"8DA4716B",
x"8DD0721D",
x"8E1A72CB",
x"8E7E736C",
x"8EF973F4",
x"8F81745B",
x"9010749C",
x"909574B0",
x"91087497",
x"915D7452",
x"919073E6",
x"919B735C",
x"918472BE",
x"9153721A",
x"91147180",
x"90D370FF",
x"909D709F",
x"907A7066",
x"906D7057",
x"90747066",
x"908A708D",
x"90A270BA",
x"90B270DC",
x"90B270EB",
x"909A70DB",
x"906C70B0",
x"902F7070",
x"8FEE702A",
x"8FBB6FEF",
x"8FA16FCF",
x"8FAC6FD9",
x"8FE37012",
x"90417075",
x"90BB70F6",
x"91407186",
x"91BF720D",
x"92217275",
x"925872AB",
x"925972A7",
x"92247266",
x"91BB71EF",
x"9128714D",
x"90737090",
x"8FA46FC5",
x"8EBB6EF6",
x"8DB46E24",
x"8C7E6D4E",
x"8B0E6C68",
x"89506B65",
x"873B6A3D",
x"84CE68E8",
x"8215676B",
x"7F2E65D0",
x"7C3E6432",
x"797962AA",
x"77106156",
x"75346055",
x"74095FBC",
x"73A35F9A",
x"74035FEE",
x"751A60B1",
x"76C661CB",
x"78E06325",
x"7B3B64A5",
x"7DAE6630",
x"801A67B4",
x"826D6926",
x"84A56A7F",
x"86C86BC4",
x"88E96CFD",
x"8B1D6E35",
x"8D796F78",
x"900E70D1",
x"92E37247",
x"95F173DC",
x"992E7592",
x"9C807761",
x"9FCC7944",
x"A2F47B30",
x"A5E07D18",
x"A8777EF0",
x"AAB280A9",
x"AC8B823C",
x"AE0E839E",
x"AF4C84C7",
x"B05B85B9",
x"B1598677",
x"B2608708",
x"B3878777",
x"B4DE87D3",
x"B66D8829",
x"B8328885",
x"BA1C88F0",
x"BC188969",
x"BE0789EC",
x"BFC78A6D",
x"C13A8ADD",
x"C2468B2A",
x"C2D88B42",
x"C2EA8B1A",
x"C2858AAE",
x"C1BC8A01",
x"C0AF8921",
x"BF888821",
x"BE708718",
x"BD948627",
x"BD168564",
x"BD1484E8",
x"BD9884C2",
x"BEA284F8",
x"C0228588",
x"C1F88663",
x"C3FE8774",
x"C60588A1",
x"C7E089CA",
x"C9658AD3",
x"CA758BA1",
x"CAFB8C21",
x"CAEF8C48",
x"CA5B8C15",
x"C9578B97",
x"C8048ADD",
x"C6888A08",
x"C5128936",
x"C3CD8888",
x"C2D8881D",
x"C2508805",
x"C23C884C",
x"C29988ED",
x"C35889D8",
x"C4598AEF",
x"C5778C13",
x"C68B8D1D",
x"C76E8DEF",
x"C8068E6F",
x"C8408E91",
x"C8188E53",
x"C7968DC3",
x"C6D38CF6",
x"C5E88C07",
x"C4F48B10",
x"C4128A29",
x"C3538967",
x"C2BD88D2",
x"C24C8869",
x"C1ED8827",
x"C1858800",
x"C0FC87E4",
x"C03587C9",
x"BF2087A2",
x"BDB78769",
x"BC028718",
x"BA1686B2",
x"B8148638",
x"B62285AC",
x"B4678514",
x"B3088473",
x"B21F83CF",
x"B1BC832D",
x"B1DE8297",
x"B2788215",
x"B36E81B0",
x"B49B8172",
x"B5D6815E",
x"B6F48178",
x"B7CC81BC",
x"B83C821C",
x"B82D828A",
x"B79882EE",
x"B6788335",
x"B4DA8346",
x"B2D18314",
x"B074828E",
x"ADD681B3",
x"AB088080",
x"A8117EFA",
x"A4ED7D25",
x"A18D7B06",
x"9DDA78A5",
x"99C075FF",
x"95287317",
x"90066FEF",
x"8A606C8A",
x"845068F6",
x"7E036544",
x"77B56194",
x"71B25E08",
x"6C495AD0",
x"67C45814",
x"645B55FE",
x"623654AD",
x"615E5432",
x"61C75489",
x"634755A3",
x"65A7575A",
x"689E5982",
x"6BEB5BE3",
x"6F445E48",
x"72776080",
x"755B6263",
x"77D663DD",
x"79E364E3",
x"7B81657C",
x"7CBE65BA",
x"7DA865B4",
x"7E506589",
x"7EC46555",
x"7F0E652F",
x"7F386528",
x"7F486549",
x"7F416594",
x"7F2A6606",
x"7F096696",
x"7EE56737",
x"7EC667DF",
x"7EB46886",
x"7EB46921",
x"7EC969AD",
x"7EF76A23",
x"7F3B6A84",
x"7F8C6ACF",
x"7FE56B04",
x"803E6B23",
x"808D6B2D",
x"80CF6B24",
x"81016B0D",
x"81246AEC",
x"813E6AC8",
x"81556AA8",
x"81726A96",
x"819B6A99",
x"81D96AB7",
x"822A6AF3",
x"828E6B4C",
x"83006BBD",
x"83746C38",
x"83E56CB4",
x"84456D21",
x"84916D70",
x"84C86D9C",
x"84F06D9D",
x"85116D78",
x"853A6D35",
x"85746CE2",
x"85D06C92",
x"86506C52",
x"86F76C31",
x"87BC6C3A",
x"88916C6B",
x"89626CBF",
x"8A1B6D30",
x"8AAA6DAB",
x"8B016E27",
x"8B1F6E97",
x"8B096EF5",
x"8ACE6F44",
x"8A846F86",
x"8A466FC7",
x"8A2C7013",
x"8A4C7075",
x"8AAF70F2",
x"8B5A718D",
x"8C467240",
x"8D6072FE",
x"8E9173B7",
x"8FC17458",
x"90D374D1",
x"91B27515",
x"924C7517",
x"929874DA",
x"9291745E",
x"923C73AF",
x"919D72D7",
x"90BF71E4",
x"8FAC70E2",
x"8E706FDB",
x"8D116ED5",
x"8B9B6DD5",
x"8A156CD9",
x"88876BE3",
x"86F96AF2",
x"85766A09",
x"840A6928",
x"82BF6856",
x"81A5679D",
x"80C96701",
x"803B668E",
x"8003664B",
x"802A663B",
x"80AF6660",
x"819066BB",
x"82BE6744",
x"842567F3",
x"85A868BA",
x"8728698C",
x"88816A5B",
x"89956B17",
x"8A496BB4",
x"8A8B6C27",
x"8A586C6B",
x"89B76C7A",
x"88B96C57",
x"877C6C02",
x"86186B82",
x"84A86ADE",
x"833F6A19",
x"81E06938",
x"8080683E",
x"7F0A6728",
x"7D5B65F3",
x"7B52649D",
x"78D1631F",
x"75C5617D",
x"72315FB9",
x"6E2B5DDF",
x"69E55BFE",
x"659C5A30",
x"619D588F",
x"5E375735",
x"5BAE563C",
x"5A3A55B8",
x"59F555B2",
x"5AE4562C",
x"5CEC571E",
x"5FDF5874",
x"63825A18",
x"678C5BED",
x"6BBD5DDC",
x"6FDB5FCB",
x"73B861AB",
x"773B6373",
x"7A586521",
x"7D0B66B8",
x"7F60683B",
x"816369AD",
x"831E6B11",
x"849A6C65",
x"85DB6D9E",
x"86E36EB7",
x"87B16FA1",
x"88467051",
x"88A270BE",
x"88CC70E6",
x"88CC70CB",
x"88AE7073",
x"887D6FEE",
x"88466F47",
x"88146E8F",
x"87EA6DD7",
x"87CB6D28",
x"87B26C8F",
x"879B6C0A",
x"877D6B9E",
x"874F6B48",
x"870A6B02",
x"86A76AC5",
x"86206A8D",
x"85746A55",
x"84A46A1A",
x"83AE69D8",
x"82956990",
x"815F6945",
x"801168F9",
x"7EB768B1",
x"7D596872",
x"7C0A6842",
x"7AD86827",
x"79D36823",
x"790D6837",
x"788D6862",
x"7859689E",
x"787368E6",
x"78D26931",
x"79686975",
x"7A2369A8",
x"7AEC69C8",
x"7BAF69D1",
x"7C5C69C2",
x"7CE269A6",
x"7D3E6982",
x"7D6F6962",
x"7D7A694E",
x"7D6F6951",
x"7D55696B",
x"7D3B699D",
x"7D2769DF",
x"7D196A26",
x"7D0E6A65",
x"7CFF6A8A",
x"7CDC6A8F",
x"7CA06A66",
x"7C416A13",
x"7BC5699A",
x"7B38690C",
x"7AB16879",
x"7A4C67FC",
x"7A3167AE",
x"7A8067A4",
x"7B5867F2",
x"7CC868A0",
x"7ED569B1",
x"81706B20",
x"847C6CDB",
x"87CD6ECF",
x"8B3870E2",
x"8E8872FC",
x"91977501",
x"944376DB",
x"96817878",
x"984C79CD",
x"99B27ACE",
x"9AC87B7C",
x"9BA27BD9",
x"9C597BE8",
x"9CFA7BB2",
x"9D8A7B40",
x"9E037A9C",
x"9E5A79D1",
x"9E8078EA",
x"9E6477F2",
x"9DFE76F4",
x"9D4B75F5",
x"9C4F74FE",
x"9B1E7412",
x"99CD7336",
x"98797268",
x"973B71AA",
x"962870FE",
x"95507064",
x"94B96FDE",
x"94636F70",
x"94406F21",
x"94406EF3",
x"944D6EE8",
x"944C6EFE",
x"94246F2E",
x"93B96F6C",
x"92F66FA4",
x"91C26FC1",
x"900E6FA7",
x"8DCC6F41",
x"8AFA6E7C",
x"879E6D4B",
x"83C86BB2",
x"7F9769BF",
x"7B32678A",
x"76CC6535",
x"729A62EA",
x"6ED460D0",
x"6BA85F0E",
x"69425DBD",
x"67B85CEE",
x"67135C9F",
x"674A5CC8",
x"68405D4F",
x"69D45E1A",
x"6BD75F08",
x"6E1B6003",
x"707760F0",
x"72C761C6",
x"74F26280",
x"76EB6324",
x"78AE63B9",
x"7A3E644E",
x"7BA764E9",
x"7CF26595",
x"7E276650",
x"7F4F671B",
x"806C67EC",
x"817D68B8",
x"82816977",
x"83726A20",
x"844F6AAB",
x"85146B1A",
x"85C56B70",
x"865F6BB2",
x"86E76BE9",
x"875F6C1A",
x"87C56C4B",
x"88176C7F",
x"88526CB1",
x"886F6CDF",
x"88696D03",
x"88396D14",
x"87E06D10",
x"87606CF3",
x"86C16CBD",
x"86116C70",
x"855F6C16",
x"84BE6BB4",
x"84416B57",
x"83F66B06",
x"83E66AC9",
x"84146AA6",
x"847A6A9C",
x"85106AAA",
x"85C26ACC",
x"867E6AFD",
x"87326B34",
x"87CD6B6B",
x"88456B9D",
x"88956BC7",
x"88C26BE8",
x"88D66C03",
x"88E06C1A",
x"88F66C37",
x"89256C5F",
x"89806C9A",
x"8A116CEF",
x"8ADA6D62",
x"8BD86DF5",
x"8CFB6EA7",
x"8E366F73",
x"8F727052",
x"9094713A",
x"918D721D",
x"924972EF",
x"92BF73A3",
x"92EF742D",
x"92DC7486",
x"929474AC",
x"9229749C",
x"91AE745E",
x"913873FB",
x"90D87382",
x"909A7300",
x"90847289",
x"90957227",
x"90C871E6",
x"910B71CB",
x"915371D2",
x"918A71F8",
x"91A17230",
x"9188726A",
x"91387296",
x"90A972A9",
x"8FE07296",
x"8EE4725A",
x"8DBF71F2",
x"8C847169",
x"8B4570C7",
x"8A137016",
x"88FD6F66",
x"88146EBF",
x"875F6E2A",
x"86E26DA9",
x"869A6D3B",
x"86806CE1",
x"86886C96",
x"86A76C58",
x"86CC6C26",
x"86E76BFD",
x"86F16BE3",
x"86E06BD5",
x"86AE6BD5",
x"865D6BDE",
x"85F06BEB",
x"856A6BF3",
x"84D26BEF",
x"842C6BD4",
x"83806B9A",
x"82CE6B3F",
x"82176AC4",
x"815B6A2E",
x"80976987",
x"7FC668D8",
x"7EE3682A",
x"7DE36781",
x"7CBF66E0",
x"7B6C6641",
x"79E06598",
x"781764DC",
x"760F6400",
x"73C862FD",
x"715161D3",
x"6EBB6087",
x"6C205F29",
x"69A15DCF",
x"67605C90",
x"65825B84",
x"64245AC0",
x"635C5A52",
x"633A5A3C",
x"63BA5A78",
x"64D15AFB",
x"66685BAF",
x"68605C82",
x"6A975D5F",
x"6CEE5E38",
x"6F455F04",
x"71895FC3",
x"73AB607A",
x"75A86132",
x"778161F7",
x"794162D0",
x"7AED63C4",
x"7C9364D5",
x"7E3565FF",
x"7FD8673A",
x"8179687C",
x"830E69B5",
x"84906ADC",
x"85F16BE6",
x"87276CCA",
x"88276D82",
x"88EF6E0D",
x"897E6E6E",
x"89DA6EA6",
x"8A0E6EBD",
x"8A286EB7",
x"8A356E9E",
x"8A456E7A",
x"8A666E54",
x"8A9F6E30",
x"8AF36E16",
x"8B606E0A",
x"8BDF6E10",
x"8C606E27",
x"8CD86E4E",
x"8D356E82",
x"8D6F6EBD",
x"8D7B6EFA",
x"8D5D6F38",
x"8D156F6F",
x"8CAF6F9F",
x"8C3B6FC3",
x"8BC56FDF",
x"8B5F6FF2",
x"8B146FFE",
x"8AE97003",
x"8AE07003",
x"8AF47000",
x"8B1B6FFA",
x"8B4B6FF0",
x"8B736FE1",
x"8B896FCD",
x"8B816FB3",
x"8B566F92",
x"8B076F6B",
x"8A986F3B",
x"8A106F08",
x"897D6ED1",
x"88EA6E9A",
x"886A6E68",
x"88066E3E",
x"87CB6E21",
x"87C16E16",
x"87E76E1E",
x"883C6E3E",
x"88B96E73",
x"89526EBB",
x"89F96F10",
x"8A9D6F6C",
x"8B2F6FC7",
x"8BA57016",
x"8BF67054",
x"8C1E7079",
x"8C217085",
x"8C067075",
x"8BD3704E",
x"8B987017",
x"8B636FD9",
x"8B3C6F9F",
x"8B316F70",
x"8B456F58",
x"8B7B6F5C",
x"8BD56F7E",
x"8C466FBD",
x"8CC97010",
x"8D4F706F",
x"8DC870CB",
x"8E227114",
x"8E4F713E",
x"8E42713D",
x"8DF47106",
x"8D65709A",
x"8C9D7000",
x"8BAB6F47",
x"8AA86E7F",
x"89AF6DC2",
x"88DC6D27",
x"88496CC2",
x"88086CA6",
x"88216CD2",
x"88916D48",
x"89486DF8",
x"8A2E6ECD",
x"8B256FAB",
x"8C13707A",
x"8CDC7123",
x"8D6F7193",
x"8DC671C4",
x"8DE371B7",
x"8DCF7175",
x"8D94710C",
x"8D3E708F",
x"8CCD7009",
x"8C3E6F83",
x"8B7A6EFE",
x"8A6C6E70",
x"88F26DCD",
x"86F06CFF",
x"84536BF0",
x"81136A96",
x"7D3768E6",
x"78DF66E6",
x"743564A3",
x"6F756235",
x"6AE15FBE",
x"66B85D60",
x"63365B3D",
x"60835974",
x"5EBD5817",
x"5DEC572E",
x"5E0556B8",
x"5EEE56AB",
x"608356F7",
x"629C578A",
x"65065850",
x"679A593C",
x"6A315A43",
x"6CAD5B60",
x"6EF65C90",
x"71015DD2",
x"72C95F25",
x"744F6081",
x"759E61E0",
x"76C46332",
x"77CF646A",
x"78D56577",
x"79E5664E",
x"7B1066E8",
x"7C636745",
x"7DE5676D",
x"7F966772",
x"81706765",
x"83696760",
x"85706777",
x"877067BB",
x"89506832",
x"8AFA68DC",
x"8C5A69AE",
x"8D606A99",
x"8E016B82",
x"8E3B6C55",
x"8E106CFD",
x"8D8E6D69",
x"8CC36D93",
x"8BC56D7A",
x"8AA86D26",
x"89806CA6",
x"885F6C0A",
x"87536B65",
x"86666AC8",
x"859A6A41",
x"84ED69D5",
x"845D6989",
x"83E5695B",
x"837D6947",
x"83216947",
x"82D06955",
x"828D696C",
x"8259698A",
x"823E69AD",
x"823F69D2",
x"826569FC",
x"82B26A2B",
x"83276A5B",
x"83BF6A8C",
x"84766ABA",
x"85416AE1",
x"86166AFC",
x"86E96B0A",
x"87B16B0A",
x"88666B00",
x"89066AED",
x"89906ADB",
x"8A066ACE",
x"8A6F6AD1",
x"8AD06AE8",
x"8B346B19",
x"8B9E6B65",
x"8C186BCB",
x"8CA46C47",
x"8D466CD4",
x"8DFC6D6B",
x"8EC56E05",
x"8F9D6E9D",
x"907E6F31",
x"91626FC0",
x"92407045",
x"931270C5",
x"93CF7140",
x"946D71B5",
x"94E67226",
x"9535728F",
x"955572F1",
x"95437347",
x"9503738D",
x"949273C1",
x"93FA73DC",
x"933E73DC",
x"926473BD",
x"9179737C",
x"90817317",
x"8F877290",
x"8E9271E6",
x"8DAE7120",
x"8CE07047",
x"8C326F65",
x"8BAA6E8A",
x"8B4C6DC5",
x"8B186D27",
x"8B106CBD",
x"8B2A6C8D",
x"8B5A6C9E",
x"8B976CEC",
x"8BCC6D6B",
x"8BEA6E08",
x"8BE26EAE",
x"8BA86F47",
x"8B366FBA",
x"8A896FF3",
x"89A46FE9",
x"888D6F93",
x"874D6EF6",
x"85EC6E17",
x"846D6D06",
x"82D56BCF",
x"811E6A82",
x"7F456928",
x"7D4167C9",
x"7B0E6668",
x"78A86500",
x"7614638D",
x"735C620A",
x"70906072",
x"6DC55EC3",
x"6B195D04",
x"68A35B3F",
x"667A5981",
x"64B457E0",
x"6358566E",
x"62695542",
x"61E25468",
x"61B553EE",
x"61D553D4",
x"62315418",
x"62B854AC",
x"63615581",
x"64235682",
x"64FA579B",
x"65E658BA",
x"66E659D3",
x"67FA5ADA",
x"691E5BCD",
x"6A4E5CAC",
x"6B805D7A",
x"6CA65E3C",
x"6DB55EF3",
x"6EA05F9F",
x"6F5E603F",
x"6FE660CB",
x"7038613B",
x"70586187",
x"704E61AB",
x"702661A5",
x"6FED6177",
x"6FB4612E",
x"6F8760D5",
x"6F72607D",
x"6F7D6038",
x"6FAB6014",
x"6FFF6018",
x"7072604B",
x"70FF60A4",
x"71986118",
x"7238619A",
x"72D16214",
x"73586277",
x"73CB62B7",
x"742462CB",
x"746362B4",
x"74906276",
x"74AB621E",
x"74C161B7",
x"74D2614F",
x"74E660F3",
x"74FF60AB",
x"7519607E",
x"7531606A",
x"75426070",
x"75476088",
x"753C60B1",
x"752160E2",
x"74F96115",
x"74C9614B",
x"749B617D",
x"747961AB",
x"746961D2",
x"747461F3",
x"749A620B",
x"74D6621D",
x"75246227",
x"75736229",
x"75BB6225",
x"75EC621E",
x"75FD6215",
x"75EA620A",
x"75B261FD",
x"755961ED",
x"74EA61DC",
x"747261C6",
x"73F961AD",
x"738C618E",
x"73356170",
x"72F76153",
x"72D6613C",
x"72CF6131",
x"72DF6134",
x"73006143",
x"732D6162",
x"73606184",
x"739361A5",
x"73C161BC",
x"73E261BE",
x"73EF61A5",
x"73E0616F",
x"73B2611D",
x"735C60B5",
x"72DB6043",
x"72315FD5",
x"71655F74",
x"707D5F2C",
x"6F8A5F06",
x"6E9E5EFE",
x"6DC95F15",
x"6D205F42",
x"6CAA5F78",
x"6C735FB1",
x"6C785FDD",
x"6CB35FF9",
x"6D135FFD",
x"6D865FE7",
x"6DF55FB9",
x"6E475F76",
x"6E6C5F1F",
x"6E545EB7",
x"6DF85E3F",
x"6D595DBC",
x"6C835D2F",
x"6B845C9A",
x"6A6F5C04",
x"695B5B70",
x"685B5AE6",
x"67805A69",
x"66D559FD",
x"665C599F",
x"660F594C",
x"65DC58F7",
x"65B15892",
x"6570580C",
x"64FF5756",
x"64425664",
x"63265532",
x"61A153C4",
x"5FB7522F",
x"5D7C5089",
x"5B0F4EF8",
x"589F4D9F",
x"565D4CA2",
x"54804C1F",
x"53384C29",
x"52AA4CC4",
x"52E84DE8",
x"53F34F7C",
x"55B75161",
x"5810536D",
x"5ACC5577",
x"5DB5575D",
x"60945904",
x"633B5A5C",
x"65895B60",
x"67695C18",
x"68DB5C91",
x"69E95CDC",
x"6AA45D0D",
x"6B285D2F",
x"6B8C5D4F",
x"6BE35D6E",
x"6C3F5D90",
x"6CA75DAE",
x"6D205DC5",
x"6DA55DD0",
x"6E375DD2",
x"6ECC5DCB",
x"6F625DC2",
x"6FF55DC1",
x"707F5DCD",
x"70FF5DEE",
x"716F5E24",
x"71CC5E6C",
x"72105EBF",
x"72375F14",
x"723E5F5C",
x"72245F91",
x"71EF5FAB",
x"71A75FA8",
x"71565F8B",
x"710A5F5C",
x"70CF5F25",
x"70AE5EF3",
x"70AD5ECF",
x"70CC5EC1",
x"71045EC9",
x"714F5EEC",
x"719D5F22",
x"71E55F66",
x"721C5FB2",
x"723D6000",
x"724B604C",
x"724B6097",
x"724960E2",
x"7251612E",
x"726D617E",
x"72A861D0",
x"73026225",
x"73766274",
x"73FA62B7",
x"747F62E4",
x"74ED62F3",
x"753862DD",
x"754C629E",
x"75236239",
x"74BB61B4",
x"741D611B",
x"7358607E",
x"72835FEE",
x"71B75F7C",
x"710A5F33",
x"70915F1E",
x"70595F42",
x"70655F9B",
x"70B1601F",
x"712E60C2",
x"71CC6173",
x"7272621D",
x"730C62AE",
x"73846318",
x"73D2634C",
x"73EC6348",
x"73D56309",
x"73966298",
x"733B6201",
x"72D66156",
x"727660A9",
x"722B6010",
x"71FD5F98",
x"71F25F53",
x"72045F45",
x"722E5F72",
x"72615FCF",
x"728A6055",
x"729D60F2",
x"728A6194",
x"72476229",
x"71D162A4",
x"713062F4",
x"70706318",
x"6FA7630A",
x"6EED62D0",
x"6E5F6270",
x"6E1661F6",
x"6E25616C",
x"6E9660E2",
x"6F696060",
x"70945FF6",
x"72025FA8",
x"73935F7D",
x"75285F77",
x"76A15F95",
x"77DD5FD2",
x"78C86024",
x"794E6081",
x"796660DC",
x"79136125",
x"7855614F",
x"7738614F",
x"75C6611D",
x"740D60B4",
x"72186014",
x"6FF75F43",
x"6DBB5E4D",
x"6B765D3D",
x"693C5C24",
x"67295B12",
x"65555A17",
x"63DC5945",
x"62D458A6",
x"624C5849",
x"624E5833",
x"62D5586A",
x"63D958EE",
x"654459B9",
x"66FA5AC2",
x"68E25BFA",
x"6AE15D4F",
x"6CDC5EAE",
x"6ECB6001",
x"70A76139",
x"72726248",
x"74386327",
x"760A63DC",
x"77F76470",
x"7A1164F6",
x"7C606586",
x"7EE96638",
x"81A86723",
x"848E6859",
x"878D69E1",
x"8A8B6BB5",
x"8D716DCB",
x"90297008",
x"929F724D",
x"94C57478",
x"96927668",
x"98087803",
x"992E7939",
x"9A0D7A03",
x"9AB57A6B",
x"9B3B7A7F",
x"9BAE7A5B",
x"9C1C7A1F",
x"9C9279E5",
x"9D1879CA",
x"9DAF79DE",
x"9E507A28",
x"9EF77AA6",
x"9F997B4D",
x"A02B7C09",
x"A0A47CC4",
x"A0FB7D6A",
x"A1307DE5",
x"A1457E2A",
x"A13B7E36",
x"A11F7E09",
x"A0FA7DAF",
x"A0D67D35",
x"A0BF7CAD",
x"A0B97C2A",
x"A0CC7BBA",
x"A0F47B6B",
x"A1347B40",
x"A1807B3A",
x"A1D07B57",
x"A21B7B89",
x"A2527BC6",
x"A2647BFC",
x"A2487C1E",
x"A1EE7C18",
x"A14D7BE1",
x"A0617B72",
x"9F297AC6",
x"9DAC79E3",
x"9BF878D1",
x"9A2277A2",
x"98427665",
x"96707534",
x"94C8741F",
x"935A7336",
x"92357280",
x"915D7202",
x"90CB71B4",
x"9070718A",
x"90397175",
x"90117161",
x"8FE47140",
x"8FA87108",
x"8F5670B7",
x"8EF17055",
x"8E876FEE",
x"8E276F93",
x"8DE66F59",
x"8DD36F52",
x"8DF96F8D",
x"8E5C700A",
x"8EF670CA",
x"8FB771B9",
x"908872C5",
x"915273D2",
x"91FE74C7",
x"9276758B",
x"92AF760B",
x"92A47641",
x"925A762D",
x"91DF75DC",
x"91437562",
x"90A274D7",
x"90137454",
x"8FA873F4",
x"8F7673C6",
x"8F8373D2",
x"8FD27419",
x"9058748F",
x"91017520",
x"91B875B0",
x"925A7626",
x"92C97665",
x"92E7765A",
x"929E75F6",
x"91E0753B",
x"90AF7431",
x"8F1A72EB",
x"8D397180",
x"8B31700D",
x"89276EAD",
x"873E6D75",
x"85936C6D",
x"842C6B9A",
x"83076AF0",
x"82076A5B",
x"810169BE",
x"7FC168FA",
x"7E0E67F3",
x"7BBB6693",
x"78A464CB",
x"74C2629A",
x"702A6011",
x"6B095D49",
x"65A95A67",
x"605F5798",
x"5B8F550B",
x"578F52E7",
x"54AA5150",
x"530F505B",
x"52D05012",
x"53DB506E",
x"5606515B",
x"590D52C0",
x"5C9D5475",
x"60655659",
x"64165846",
x"67735A21",
x"6A545BD2",
x"6CA75D4B",
x"6E705E87",
x"6FC45F87",
x"70C16052",
x"718C60F3",
x"72476172",
x"730A61D8",
x"73E6622E",
x"74E2627A",
x"75F762BF",
x"771A6300",
x"783A633E",
x"7948637F",
x"7A3963C2",
x"7B04640E",
x"7BA86466",
x"7C2564CF",
x"7C846548",
x"7CCC65D2",
x"7D066669",
x"7D386707",
x"7D6867A5",
x"7D956838",
x"7DC568B8",
x"7DF3691E",
x"7E1E6963",
x"7E446983",
x"7E636980",
x"7E7C6959",
x"7E8B6914",
x"7E9468B5",
x"7E916841",
x"7E8767BC",
x"7E736730",
x"7E58669D",
x"7E3A660E",
x"7E1B6589",
x"7E016518",
x"7DF564C4",
x"7DFC6497",
x"7E18649B",
x"7E5264D5",
x"7EA76548",
x"7F1365EF",
x"7F9166C2",
x"801A67B1",
x"80A068AA",
x"811B6999",
x"81816A65",
x"81CB6AFF",
x"81F46B59",
x"81FE6B6D",
x"81EA6B3F",
x"81BE6AD8",
x"81816A47",
x"813B69A0",
x"80F368F7",
x"80B16862",
x"807C67ED",
x"805867A1",
x"80456781",
x"80456787",
x"805567AD",
x"806C67E0",
x"80846819",
x"80976846",
x"8097685F",
x"807E685E",
x"8049683F",
x"7FF66807",
x"7F8467BA",
x"7EFC675E",
x"7E6766FC",
x"7DD2669B",
x"7D466644",
x"7CCF65F5",
x"7C6F65B1",
x"7C256577",
x"7BEF6545",
x"7BBF6517",
x"7B8A64E9",
x"7B4164BA",
x"7AD66487",
x"7A456455",
x"798A6423",
x"78A863F3",
x"77AB63C9",
x"769E63AA",
x"75946390",
x"749B637C",
x"73C16369",
x"7311634F",
x"72906328",
x"723D62EC",
x"72166293",
x"7211621B",
x"722A6187",
x"725160D9",
x"727F601A",
x"72A85F56",
x"72C45E9B",
x"72C95DF6",
x"72B05D70",
x"72705D10",
x"72065CD5",
x"71695CBB",
x"70975CB8",
x"6F8D5CB9",
x"6E4A5CAE",
x"6CCF5C82",
x"6B1D5C26",
x"69385B8E",
x"67275AB5",
x"64EE599E",
x"62975852",
x"603056E3",
x"5DC5556A",
x"5B6E53FD",
x"594052B9",
x"575851B5",
x"55D15101",
x"54C550AC",
x"544D50B6",
x"5473511B",
x"553D51CD",
x"56A252BD",
x"588953D4",
x"5AD454FD",
x"5D585621",
x"5FEB5732",
x"625E5824",
x"648D58F1",
x"665F599C",
x"67C55A28",
x"68BE5A9E",
x"69585B05",
x"69A65B6A",
x"69C75BCF",
x"69D55C36",
x"69EB5CA4",
x"6A1D5D10",
x"6A735D78",
x"6AF35DD6",
x"6B945E25",
x"6C4B5E62",
x"6D095E8E",
x"6DBD5EAE",
x"6E585EC3",
x"6ECF5ED7",
x"6F1B5EF0",
x"6F3E5F14",
x"6F3C5F45",
x"6F1D5F87",
x"6EEF5FD8",
x"6EBF6032",
x"6E9D6094",
x"6E9660F7",
x"6EB46156",
x"6F0061AF",
x"6F7C6200",
x"70266248",
x"70F96289",
x"71E962C2",
x"72E962F9",
x"73EC632D",
x"74E0635D",
x"75BA638B",
x"766F63B7",
x"76FA63DF",
x"775E6404",
x"779D6425",
x"77BF6444",
x"77D36462",
x"77E66480",
x"780664A0",
x"783E64C2",
x"789764E6",
x"7916650A",
x"79BE652E",
x"7A8C654E",
x"7B796568",
x"7C7F657D",
x"7D91658E",
x"7EA865A0",
x"7FB765B5",
x"80B565D2",
x"819B65FD",
x"82656638",
x"83106684",
x"839B66DF",
x"840A6746",
x"846267B2",
x"84A4681B",
x"84D6687A",
x"84F768C9",
x"850A6900",
x"8509691B",
x"84EF691B",
x"84B568FF",
x"845968C7",
x"83D36877",
x"83256816",
x"825267A7",
x"81606735",
x"805F66C6",
x"7F596668",
x"7E626620",
x"7D8465FA",
x"7CCB65FF",
x"7C3B6630",
x"7BD5668E",
x"7B936713",
x"7B6967B2",
x"7B4E685B",
x"7B3568FA",
x"7B18697C",
x"7AF369CE",
x"7AC469E1",
x"7A8E69B1",
x"7A58693E",
x"7A2A6890",
x"7A0467B5",
x"79ED66C4",
x"79DD65CF",
x"79D164EA",
x"79BC6425",
x"7996638D",
x"79536325",
x"78F062ED",
x"786B62DF",
x"77C862F3",
x"770E631B",
x"764B634C",
x"7589637A",
x"74CF6397",
x"74216397",
x"737A6372",
x"72D3631D",
x"721C6294",
x"714461D5",
x"703E60E0",
x"6F045FC1",
x"6D965E80",
x"6BFC5D33",
x"6A4E5BF0",
x"68A65ACF",
x"672459E4",
x"65E65945",
x"650958FD",
x"649A590F",
x"64A15975",
x"65175A21",
x"65E85AF8",
x"66F95BE4",
x"682D5CCB",
x"69685D94",
x"6A8F5E31",
x"6B935E9D",
x"6C6C5ED6",
x"6D1E5EEA",
x"6DB35EE7",
x"6E3A5EE0",
x"6EC55EE6",
x"6F655F06",
x"70245F4B",
x"710C5FB7",
x"721C6048",
x"734F60F7",
x"74A161BC",
x"7606628E",
x"77726363",
x"78DB6437",
x"7A326503",
x"7B7265C6",
x"7C8D667F",
x"7D7C6728",
x"7E3467C4",
x"7EB26849",
x"7EF168B5",
x"7EF56903",
x"7EBE692E",
x"7E5D693B",
x"7DE3692A",
x"7D666907",
x"7CFF68E1",
x"7CC668C2",
x"7CD468BE",
x"7D3868E1",
x"7DFA6931",
x"7F1D69B1",
x"80936A5B",
x"824C6B20",
x"842F6BEF",
x"86246CB3",
x"880D6D59",
x"89D36DD2",
x"8B656E14",
x"8CB46E1D",
x"8DBB6DF5",
x"8E796DA7",
x"8EF36D44",
x"8F326CDE",
x"8F3F6C84",
x"8F256C44",
x"8EEC6C20",
x"8E9B6C19",
x"8E396C27",
x"8DCC6C42",
x"8D566C5E",
x"8CDC6C6F",
x"8C636C6D",
x"8BF06C59",
x"8B8A6C30",
x"8B356BFA",
x"8AF96BBE",
x"8AD86B86",
x"8AD26B59",
x"8AE46B3F",
x"8B0B6B3B",
x"8B3C6B4C",
x"8B6F6B70",
x"8B976BA6",
x"8BAC6BE6",
x"8BAA6C33",
x"8B8E6C86",
x"8B5D6CE2",
x"8B226D48",
x"8AE66DB8",
x"8AB66E30",
x"8A9F6EB0",
x"8AAB6F31",
x"8ADA6FAE",
x"8B2A701F",
x"8B90707C",
x"8BFD70BD",
x"8C6370DC",
x"8CAF70D8",
x"8CD370B1",
x"8CC8706B",
x"8C86700A",
x"8C146F97",
x"8B796F1A",
x"8ABF6E99",
x"89F66E1C",
x"892B6DA6",
x"88676D3E",
x"87B56CE9",
x"871B6CA7",
x"869D6C7D",
x"863C6C6D",
x"85FC6C76",
x"85DB6C96",
x"85DC6CCA",
x"85FE6D0A",
x"863F6D51",
x"869B6D8F",
x"87086DBD",
x"87806DCE",
x"87F26DBB",
x"88506D80",
x"888E6D1D",
x"889F6C94",
x"88796BF0",
x"88136B3A",
x"87696A7A",
x"867669B8",
x"853468F6",
x"839D6830",
x"81A8675E",
x"7F4C666D",
x"7C7F654F",
x"793563F2",
x"75706248",
x"7134604B",
x"6C905DFE",
x"67A45B73",
x"629658C3",
x"5D995612",
x"58E55388",
x"54B35150",
x"51364F8F",
x"4E974E60",
x"4CF54DD1",
x"4C554DE4",
x"4CB44E89",
x"4DF54FA6",
x"4FF35116",
x"527B52B2",
x"55555453",
x"584F55D6",
x"5B365724",
x"5DE2582F",
x"603B58F8",
x"6234598A",
x"63CE59F1",
x"65145A46",
x"661A5A9E",
x"66F95B08",
x"67C75B90",
x"68995C38",
x"697B5CF8",
x"6A735DC6",
x"6B7A5E8E",
x"6C875F3C",
x"6D865FBE",
x"6E636007",
x"6F106013",
x"6F7C5FDF",
x"6FA35F76",
x"6F8A5EE9",
x"6F3C5E48",
x"6ECF5DA8",
x"6E585D1C",
x"6DF05CB3",
x"6DAD5C74",
x"6DA05C61",
x"6DD25C7B",
x"6E415CBB",
x"6EE85D17",
x"6FB75D8A",
x"709B5E0D",
x"71835E9D",
x"725F5F38",
x"73215FDD",
x"73C26091",
x"74416150",
x"74A5621B",
x"74F462ED",
x"753C63BE",
x"75876484",
x"75DF6538",
x"764865CC",
x"76C6663A",
x"7755667A",
x"77EF668B",
x"788A6670",
x"791B662E",
x"799865CE",
x"79F66559",
x"7A2D64DC",
x"7A37645F",
x"7A1163EA",
x"79BF6386",
x"79426335",
x"78A162F6",
x"77E362C6",
x"771362A2",
x"76386284",
x"755F6262",
x"748E6235",
x"73CF61F9",
x"732761A8",
x"729A6142",
x"722860C9",
x"71D16042",
x"718A5FB3",
x"714E5F28",
x"71135EA7",
x"70CF5E3B",
x"707A5DE9",
x"700D5DB6",
x"6F875DA5",
x"6EEB5DB6",
x"6E3E5DE2",
x"6D8A5E25",
x"6CDB5E74",
x"6C3B5EC8",
x"6BB45F14",
x"6B4C5F4D",
x"6B075F6D",
x"6ADF5F67",
x"6AD25F3B",
x"6AD55EE3",
x"6AE25E66",
x"6AF05DC9",
x"6AFC5D1C",
x"6B065C6D",
x"6B115BCF",
x"6B265B52",
x"6B495B0A",
x"6B865B00",
x"6BE35B3B",
x"6C625BB9",
x"6D005C74",
x"6DB75D5A",
x"6E7A5E5C",
x"6F3E5F62",
x"6FF3605A",
x"70906132",
x"710A61DD",
x"715F6256",
x"7191629B",
x"71A662B1",
x"71A4629D",
x"71946268",
x"7177621A",
x"715261BC",
x"711B6152",
x"70C860DD",
x"7046605C",
x"6F865FCC",
x"6E725F28",
x"6CF95E6C",
x"6B175D94",
x"68C85C9C",
x"661A5B87",
x"63215A57",
x"5FFF5915",
x"5CD957CC",
x"59DC568A",
x"5737555D",
x"55135457",
x"53925389",
x"52CE5302",
x"52D452CC",
x"53A452E8",
x"5531535A",
x"57655416",
x"5A1C5514",
x"5D2E5640",
x"6072578A",
x"63BB58DC",
x"66E25A26",
x"69C85B5C",
x"6C525C73",
x"6E725D64",
x"701E5E32",
x"715C5EDC",
x"72325F66",
x"72AE5FD6",
x"72E0602F",
x"72D96076",
x"72A860AD",
x"725C60D2",
x"720060EA",
x"719C60F6",
x"713760F6",
x"70D460F0",
x"707660E9",
x"702360E4",
x"6FD960EA",
x"6FA06100",
x"6F796129",
x"6F6B616C",
x"6F7C61C8",
x"6FAE623B",
x"700962C5",
x"708F635F",
x"713C6403",
x"721364A8",
x"730C6548",
x"741B65D6",
x"753B664E",
x"765B66A5",
x"777366DB",
x"787766EC",
x"796366DC",
x"7A3766B2",
x"7AF36679",
x"7BA1663B",
x"7C4C6609",
x"7D0165ED",
x"7DCC65F5",
x"7EB46624",
x"7FBF667F",
x"80EA6700",
x"822E67A1",
x"837D6854",
x"84C9690C",
x"860169BB",
x"87146A55",
x"87F96AD5",
x"88A76B37",
x"891D6B7D",
x"895C6BAE",
x"896D6BD5",
x"89566BF8",
x"89246C20",
x"88DD6C54",
x"88876C93",
x"88276CDE",
x"87BC6D2B",
x"87466D73",
x"86C56DAD",
x"86346DCD",
x"85946DCA",
x"84E36DA3",
x"84226D52",
x"83566CDC",
x"82816C47",
x"81A86B97",
x"80D16AD9",
x"7FFF6A14",
x"7F3A6952",
x"7E866897",
x"7DE667E9",
x"7D5F674B",
x"7CF066BA",
x"7C996634",
x"7C5565B8",
x"7C1E6542",
x"7BEF64CE",
x"7BBE645C",
x"7B8463EC",
x"7B396381",
x"7ADB631F",
x"7A6562CB",
x"79DB628A",
x"79426262",
x"78A06252",
x"77FC625C",
x"775B627D",
x"76C462AB",
x"763562DD",
x"75B1630B",
x"75326327",
x"74B46327",
x"742E6304",
x"739B62B8",
x"72FA6246",
x"724861B1",
x"71896101",
x"70BE6041",
x"6FF05F7D",
x"6F285EC3",
x"6E6A5E1B",
x"6DBD5D8E",
x"6D1E5D1F",
x"6C905CCB",
x"6C095C8D",
x"6B7F5C5C",
x"6AE85C2C",
x"6A355BF3",
x"695F5BA5",
x"685E5B3D",
x"67305AB8",
x"65D95A1A",
x"6468596B",
x"62EC58BC",
x"617F581C",
x"6037579C",
x"5F31574D",
x"5E83573D",
x"5E415773",
x"5E7657F1",
x"5F2758B3",
x"604F59AE",
x"61DF5AD0",
x"63C75C08",
x"65EE5D41",
x"68385E69",
x"6A905F72",
x"6CDF6050",
x"6F146104",
x"7124618D",
x"730961F4",
x"74C46245",
x"7656628B",
x"77C962D5",
x"7921632E",
x"7A63639E",
x"7B986427",
x"7CC164CB",
x"7DE06581",
x"7EFC6646",
x"80176711",
x"813B67D9",
x"8273689A",
x"83CC6955",
x"85566A0C",
x"87246AC7",
x"89416B8D",
x"8BB56C6C",
x"8E806D6C",
x"91986E93",
x"94EA6FE2",
x"98597154",
x"9BC272DE",
x"9EFE7472",
x"A1EB75FE",
x"A46D776C",
x"A66B78B0",
x"A7E179BC",
x"A8D17A85",
x"A94F7B0E",
x"A9707B5A",
x"A95A7B77",
x"A92C7B74",
x"A90A7B63",
x"A90C7B56",
x"A9497B5B",
x"A9C67B7E",
x"AA827BC4",
x"AB767C2F",
x"AC8F7CB4",
x"ADBA7D4A",
x"AEE47DE4",
x"AFF87E72",
x"B0EB7EEA",
x"B1B67F3F",
x"B2597F75",
x"B2DC7F8F",
x"B34D7F9C",
x"B3C07FAB",
x"B4497FCF",
x"B4F7801B",
x"B5D9809B",
x"B6F48157",
x"B8438249",
x"B9BA8366",
x"BB4A8498",
x"BCD785C5",
x"BE4C86D2",
x"BF9287A8",
x"C09B8838",
x"C1618881",
x"C1EA8887",
x"C2438860",
x"C2818825",
x"C2BD87F4",
x"C30F87EA",
x"C389881B",
x"C4348895",
x"C5128956",
x"C6138A4F",
x"C7258B6A",
x"C8268C88",
x"C8F78D86",
x"C9798E43",
x"C9938EA7",
x"C9348EA2",
x"C8588E31",
x"C7068D59",
x"C5538C2F",
x"C35B8ACC",
x"C1448950",
x"BF3387DA",
x"BD508688",
x"BBBA8573",
x"BA8E84A9",
x"B9DA8435",
x"B9A28415",
x"B9DC8442",
x"BA7584AC",
x"BB50853F",
x"BC4785E9",
x"BD33868F",
x"BDEE8722",
x"BE57878D",
x"BE5487C3",
x"BDD787BE",
x"BCE08776",
x"BB7786EC",
x"B9AC8623",
x"B798851F",
x"B54D83E8",
x"B2E08282",
x"B05480F5",
x"ADAB7F45",
x"AAD47D74",
x"A7BA7B84",
x"A4457977",
x"A05A774A",
x"9BF074FF",
x"97067299",
x"91AB7017",
x"8C076D83",
x"86526AE2",
x"80CC6844",
x"7BBF65B8",
x"776F6353",
x"74136128",
x"71D55F52",
x"70C25DE0",
x"70D55CE9",
x"71F05C76",
x"73E85C91",
x"76835D39",
x"798A5E67",
x"7CCC6010",
x"801E6221",
x"836C6487",
x"86AC672B",
x"89E669FA",
x"8D2E6CE2",
x"909D6FD2",
x"944C72C1",
x"985075A6",
x"9CB5787E",
x"A17B7B43",
x"A6977DF7",
x"ABEE8096",
x"B1618322",
x"B6CD8599",
x"BC0987F9",
x"C0F28A3F",
x"C56D8C6C",
x"C9648E7A",
x"CCD0906D",
x"CFB49241",
x"D21993F8",
x"D4109590",
x"D5B09707",
x"D70C985E",
x"D833998F",
x"D9319A96",
x"DA0B9B6F",
x"DABE9C16",
x"DB419C85",
x"DB899CBB",
x"DB8C9CB8",
x"DB449C82",
x"DAAD9C1A",
x"D9D19B8D",
x"D8C09AE4",
x"D78F9A2A",
x"D65E996E",
x"D54A98B8",
x"D4719817",
x"D3EC9790",
x"D3CD972D",
x"D41696F0",
x"D4C696DF",
x"D5CB96FA",
x"D70D9741",
x"D86E97AD",
x"D9CB9837",
x"DAFE98D2",
x"DBE5996C",
x"DC6599F3",
x"DC6A9A54",
x"DBE59A79",
x"DADB9A54",
x"D95899DE",
x"D7759917",
x"D554980A",
x"D32396CC",
x"D112957A",
x"CF509434",
x"CE08931B",
x"CD58924C",
x"CD5391DB",
x"CDF691D1",
x"CF2F9227",
x"D0D492CB",
x"D2B293A3",
x"D48B9487",
x"D61D9555",
x"D73095E8",
x"D7989627",
x"D73A9602",
x"D6159576",
x"D43B9490",
x"D1DA9365",
x"CF269213",
x"CC6290B9",
x"C9D48F7C",
x"C7B08E71",
x"C6268DB1",
x"C5498D42",
x"C51C8D25",
x"C58B8D52",
x"C6758DB9",
x"C7AC8E4B",
x"C9048EF4",
x"CA548FA5",
x"CB7F9055",
x"CC7890FC",
x"CD3D9198",
x"CDDB922E",
x"CE6A92C1",
x"CEFE9353",
x"CFA793E5",
x"D0719474",
x"D15494F9",
x"D2409568",
x"D31695B5",
x"D3BA95D5",
x"D40995C1",
x"D3EE9576",
x"D35D94F8",
x"D25D9453",
x"D101939A",
x"CF6492DF",
x"CDA99234",
x"CBEB91A5",
x"CA379135",
x"C88C90DB",
x"C6D39080",
x"C4DD9004",
x"C2748F3E",
x"BF5A8E06",
x"BB578C38",
x"B64689B9",
x"B0188685",
x"A8E782A8",
x"A0E67E40",
x"98697981",
x"8FDA74A7",
x"87AF6FF5",
x"80556BAD",
x"7A2A6803",
x"7572651B",
x"724C630D",
x"70B761D6",
x"708D6166",
x"7193619F",
x"73796263",
x"75F3638D",
x"78B764FC",
x"7B8C669D",
x"7E4B685E",
x"80E56A37",
x"835A6C24",
x"85BB6E20",
x"88187023",
x"8A867220",
x"8D0D7400",
x"8FAC75AF",
x"9258770F",
x"94F9780D",
x"9773789B",
x"99A778B4",
x"9B7D786A",
x"9CE777D1",
x"9DE37712",
x"9E7A7657",
x"9EC075CB",
x"9ED67597",
x"9EDC75D2",
x"9EF17688",
x"9F3277B3",
x"9FAE793E",
x"A06D7B05",
x"A16B7CE1",
x"A29A7EA5",
x"A3E68026",
x"A538814C",
x"A6778200",
x"A78F8239",
x"A87181FE",
x"A911815D",
x"A96E806A",
x"A9887F3F",
x"A9667DF7",
x"A90C7CA6",
x"A8887B64",
x"A7E37A40",
x"A7247947",
x"A6567881",
x"A58177F1",
x"A4AC7798",
x"A3E37772",
x"A32C777B",
x"A29277A6",
x"A21E77EC",
x"A1D57843",
x"A1BB789F",
x"A1CD78F7",
x"A2087947",
x"A260798C",
x"A2C579C6",
x"A32679F7",
x"A3737A22",
x"A39C7A4A",
x"A39B7A71",
x"A36B7A98",
x"A3187ABE",
x"A2B37AE4",
x"A2577B06",
x"A2227B2C",
x"A2337B58",
x"A2A87B96",
x"A3927BF2",
x"A4FB7C7C",
x"A6E07D44",
x"A9307E54",
x"ABD67FB5",
x"AEAF8167",
x"B1A18363",
x"B48E8598",
x"B76487F1",
x"BA168A55",
x"BCA08CAA",
x"BF058ED5",
x"C14990C4",
x"C36D9263",
x"C56E93AB",
x"C7479497",
x"C8E5952B",
x"CA399569",
x"CB2C955C",
x"CBB0950E",
x"CBBF948E",
x"CB5E93E8",
x"CA9D9327",
x"C99B925C",
x"C8789196",
x"C75A90DC",
x"C664903C",
x"C5AC8FB9",
x"C53C8F55",
x"C50C8F0A",
x"C5068ECC",
x"C5068E8B",
x"C4E38E36",
x"C46E8DB8",
x"C3888D01",
x"C2158C06",
x"C00F8AC2",
x"BD828939",
x"BA89877D",
x"B74F85A3",
x"B40483C7",
x"B0DD8208",
x"AE05807E",
x"AB997F3A",
x"A9A17E46",
x"A80D7D95",
x"A6B57D15",
x"A5637CA5",
x"A3CC7C18",
x"A1A57B44",
x"9EA87A01",
x"9AA5782C",
x"958175B6",
x"8F4872A1",
x"88256F02",
x"80676B00",
x"787966CF",
x"70CC62AB",
x"69DB5ED3",
x"64105B80",
x"5FBE58DF",
x"5D17570C",
x"5C245615",
x"5CCA55F3",
x"5ECE568F",
x"61DB57CC",
x"65925980",
x"69905B81",
x"6D825DA7",
x"71205FCD",
x"743F61D8",
x"76C863AF",
x"78BA6548",
x"7A246697",
x"7B21679B",
x"7BCE6858",
x"7C4568CF",
x"7C9E690C",
x"7CE86914",
x"7D2868F5",
x"7D6368B7",
x"7D956863",
x"7DBE6806",
x"7DD967A5",
x"7DE86745",
x"7DEC66EB",
x"7DE96693",
x"7DE6663F",
x"7DE665EF",
x"7DF0659E",
x"7E066552",
x"7E2B650D",
x"7E6064D8",
x"7EA764BC",
x"7F0164C5",
x"7F6F64FD",
x"7FEF6568",
x"80816609",
x"812166DC",
x"81C867D3",
x"827068E2",
x"830E69F2",
x"839A6AEF",
x"840D6BC7",
x"84656C6C",
x"84A26CDB",
x"84D26D14",
x"84FD6D23",
x"853A6D17",
x"85986D06",
x"862A6D04",
x"86F96D21",
x"880A6D6B",
x"89556DE3",
x"8AC96E8D",
x"8C4F6F5B",
x"8DCB7040",
x"8F1E712A",
x"902E720A",
x"90E672D1",
x"913C7374",
x"913473E8",
x"90D3742D",
x"90327443",
x"8F67742F",
x"8E9073F5",
x"8DC3739D",
x"8D177331",
x"8C9772B9",
x"8C49723A",
x"8C2B71C0",
x"8C32714F",
x"8C5270F4",
x"8C7670AD",
x"8C917082",
x"8C947070",
x"8C767076",
x"8C2F708D",
x"8BC070AD",
x"8B2E70CA",
x"8A7E70D7",
x"89BC70CE",
x"88F270A3",
x"882A7055",
x"876F6FE2",
x"86C86F4D",
x"86396E9C",
x"85C96DD9",
x"85746D0D",
x"853C6C45",
x"851E6B8A",
x"85146AE3",
x"851B6A59",
x"852E69F0",
x"854869AA",
x"8562698A",
x"8579698C",
x"858769B0",
x"858A69EF",
x"857B6A44",
x"855C6AA7",
x"85276B0F",
x"84DC6B70",
x"847D6BC2",
x"840A6BFA",
x"83846C10",
x"82F26BFC",
x"82566BBD",
x"81B86B52",
x"811D6AC4",
x"808D6A1A",
x"80116963",
x"7FAE68AE",
x"7F6A680A",
x"7F466786",
x"7F41672A",
x"7F5366FC",
x"7F7066F7",
x"7F866713",
x"7F7A673B",
x"7F356758",
x"7E9B6753",
x"7D936711",
x"7C0B667D",
x"79FC658B",
x"77666435",
x"745E6286",
x"7100608D",
x"6D765E67",
x"69F65C36",
x"66B45A22",
x"63E6584D",
x"61BB56DA",
x"605655E1",
x"5FCB5570",
x"601D5588",
x"613B5625",
x"6309572F",
x"655C588F",
x"68025A25",
x"6AC85BD0",
x"6D7F5D6E",
x"6FFA5EE4",
x"721D601B",
x"73D36104",
x"7519619B",
x"75F261E3",
x"767361E8",
x"76B061B8",
x"76C6616D",
x"76CF611D",
x"76E560DD",
x"771760C2",
x"777560D6",
x"77FF6121",
x"78B4619F",
x"79876248",
x"7A6D630A",
x"7B5563D5",
x"7C2F6493",
x"7CF26534",
x"7D9365AA",
x"7E1065ED",
x"7E6D65FD",
x"7EAE65E0",
x"7EDF65A1",
x"7F06654E",
x"7F2B64F7",
x"7F5564AE",
x"7F866480",
x"7FBA6474",
x"7FED6493",
x"801B64D8",
x"803C653F",
x"804C65C4",
x"80486658",
x"802F66F3",
x"80076789",
x"7FD56810",
x"7F9E6883",
x"7F6D68DE",
x"7F48691E",
x"7F326948",
x"7F32695F",
x"7F446966",
x"7F656968",
x"7F8E6965",
x"7FBA6965",
x"7FDF6966",
x"7FF76968",
x"7FFD6968",
x"7FF0695E",
x"7FCE6944",
x"7F9D6913",
x"7F6268C8",
x"7F256863",
x"7EF367E8",
x"7ED2675E",
x"7ECB66CF",
x"7EE3664C",
x"7F1D65E2",
x"7F77659B",
x"7FF26581",
x"8089659A",
x"813265E2",
x"81EA6652",
x"82A766DE",
x"835D6776",
x"8404680D",
x"848E6896",
x"84F16903",
x"85216951",
x"8515697D",
x"84C8698C",
x"84386983",
x"836A696B",
x"826A694C",
x"814E6930",
x"8028691D",
x"7F146914",
x"7E2B6919",
x"7D836926",
x"7D256935",
x"7D196944",
x"7D556949",
x"7DCB693E",
x"7E636920",
x"7F0168EB",
x"7F8C689E",
x"7FE96841",
x"800967D6",
x"7FE6676B",
x"7F816703",
x"7EE666AB",
x"7E2A666C",
x"7D5F6646",
x"7C9D663F",
x"7BF66650",
x"7B7A6672",
x"7B2E669A",
x"7B1366BB",
x"7B2166CB",
x"7B4B66C1",
x"7B836696",
x"7BB7664B",
x"7BD565E8",
x"7BCC6575",
x"7B8C64FA",
x"7B096487",
x"7A35641D",
x"790963BF",
x"777F6368",
x"75966307",
x"734F6291",
x"70B761F3",
x"6DDB6121",
x"6AD26011",
x"67BA5EC6",
x"64B55D4D",
x"61E85BBD",
x"5F755A33",
x"5D7D58D0",
x"5C1C57B3",
x"5B5E56F5",
x"5B4A56A8",
x"5BD856CA",
x"5CF85756",
x"5E8D5835",
x"6079594A",
x"62975A7A",
x"64C95BA4",
x"66F25CAE",
x"68FC5D87",
x"6AD75E28",
x"6C7F5E92",
x"6DF05ED2",
x"6F345EF1",
x"704C5F04",
x"71425F1D",
x"721C5F46",
x"72DE5F8A",
x"738A5FEE",
x"74216070",
x"74A0610A",
x"750761AF",
x"75566256",
x"758D62F2",
x"75AB6373",
x"75B463D3",
x"75AB640A",
x"75946414",
x"757363F4",
x"754963AD",
x"751D6346",
x"74EF62CE",
x"74C2624C",
x"749D61D0",
x"74836164",
x"747A6113",
x"748D60E3",
x"74BF60DA",
x"751960FA",
x"759D6143",
x"764F61B1",
x"772E6241",
x"783562E9",
x"795963A1",
x"7A906462",
x"7BCC651D",
x"7D0065C8",
x"7E20665B",
x"7F2566C9",
x"800A6713",
x"80D36732",
x"81866731",
x"822D6714",
x"82D666EB",
x"838D66C5",
x"845C66B4",
x"854866C6",
x"86506706",
x"876D6779",
x"888E681A",
x"89A468E1",
x"8A9769BE",
x"8B556A9C",
x"8BCE6B69",
x"8BF76C13",
x"8BD36C8D",
x"8B676CD1",
x"8AC66CDF",
x"8A036CBE",
x"89386C7A",
x"887E6C24",
x"87EA6BCC",
x"878B6B83",
x"876A6B52",
x"87866B42",
x"87D66B55",
x"88506B89",
x"88E26BD8",
x"897A6C3B",
x"8A0B6CA7",
x"8A896D13",
x"8AEC6D78",
x"8B326DCE",
x"8B5F6E13",
x"8B766E44",
x"8B7F6E63",
x"8B7F6E75",
x"8B7B6E7C",
x"8B746E7F",
x"8B6A6E83",
x"8B596E8D",
x"8B3C6E9E",
x"8B0E6EBA",
x"8ACB6ED9",
x"8A736EF9",
x"8A076F13",
x"898E6F20",
x"89116F17",
x"889B6EF6",
x"88376EBB",
x"87EF6E68",
x"87C86E05",
x"87C56D9A",
x"87E36D37",
x"881A6CE3",
x"885D6CAD",
x"889E6C97",
x"88CE6CA4",
x"88DD6CCE",
x"88C16D0A",
x"886D6D48",
x"87DD6D76",
x"870D6D7F",
x"85FA6D54",
x"84A46CE3",
x"830B6C2A",
x"81316B24",
x"7F1869DB",
x"7CC86859",
x"7A4866B4",
x"77A86500",
x"74FA6355",
x"725861C6",
x"6FDE6064",
x"6DA75F3C",
x"6BD15E50",
x"6A6F5D9E",
x"69915D1E",
x"693E5CC9",
x"696D5C92",
x"6A145C73",
x"6B1D5C67",
x"6C725C6E",
x"6DFA5C90",
x"6FA45CD5",
x"71625D49",
x"732E5DF8",
x"750A5EED",
x"76FF6027",
x"791361A2",
x"7B536353",
x"7DC8652A",
x"80736710",
x"835368F2",
x"86606ABE",
x"89906C66",
x"8CCF6DE8",
x"90116F41",
x"9346707F",
x"966071AB",
x"995772D8",
x"9C287415",
x"9ED2756F",
x"A15676F1",
x"A3BB789C",
x"A6057A6F",
x"A83D7C61",
x"AA647E67",
x"AC7D806E",
x"AE848268",
x"B0778443",
x"B24D85EA",
x"B3F8874D",
x"B5708860",
x"B6A28917",
x"B78A896A",
x"B81E8959",
x"B86088EA",
x"B8578829",
x"B8118729",
x"B7A38600",
x"B72B84CC",
x"B6C483A9",
x"B68C82B6",
x"B69F820C",
x"B70B81BD",
x"B7DA81D4",
x"B904824F",
x"BA7A8321",
x"BC1C8435",
x"BDC9856E",
x"BF5386A9",
x"C09387C0",
x"C1648895",
x"C1AD890E",
x"C162891D",
x"C08888BF",
x"BF358801",
x"BD8C86FD",
x"BBBC85D4",
x"B9FA84AF",
x"B87A83B5",
x"B76A830C",
x"B6EA82CF",
x"B70A830E",
x"B7C983C9",
x"B90F84F3",
x"BABC8671",
x"BC9C8821",
x"BE7F89D9",
x"C0338B6F",
x"C18F8CBF",
x"C2758DAC",
x"C2DB8E28",
x"C2C68E2F",
x"C24D8DCE",
x"C1918D1B",
x"C0B98C38",
x"BFF18B4B",
x"BF5D8A7A",
x"BF1489E7",
x"BF2289AB",
x"BF7F89CD",
x"C0168A48",
x"C0C08B05",
x"C14E8BE2",
x"C1918CB1",
x"C15D8D43",
x"C0928D70",
x"BF258D1A",
x"BD198C35",
x"BA938ACC",
x"B7C68900",
x"B4F48700",
x"B26A850D",
x"B0738366",
x"AF4A8249",
x"AF1C81DE",
x"AFF4823B",
x"B1C08359",
x"B4528514",
x"B7608736",
x"BA92897A",
x"BD8E8B94",
x"BFFC8D3F",
x"C19B8E49",
x"C2428E97",
x"C1E78E24",
x"C0A38D0B",
x"BEA88B79",
x"BC3389A5",
x"B98C87CA",
x"B6F3861B",
x"B49184B9",
x"B27783AD",
x"B09982EE",
x"AECF8254",
x"ACDD81B0",
x"AA7880C6",
x"A7637F64",
x"A3697D63",
x"9E747AAF",
x"98977754",
x"92007378",
x"8B046F55",
x"840A6B38",
x"7D866770",
x"77E26449",
x"73786200",
x"708460B5",
x"6F1D6070",
x"6F38611E",
x"70A66290",
x"73256489",
x"766866C5",
x"7A1B6904",
x"7DFC6B10",
x"81CF6CC7",
x"85736E1D",
x"88D56F1C",
x"8BF06FDC",
x"8ECB7083",
x"916F7139",
x"93E9721C",
x"963F7345",
x"987774C0",
x"9A947683",
x"9C98787C",
x"9E877A8E",
x"A0647C94",
x"A23B7E70",
x"A4118002",
x"A5EB813D",
x"A7CD8216",
x"A9B08291",
x"AB8C82BB",
x"AD5282A5",
x"AEED826A",
x"B0508223",
x"B17081E6",
x"B24581C3",
x"B2D681CA",
x"B32F8200",
x"B3618261",
x"B38282E8",
x"B3A3838A",
x"B3D28436",
x"B41784E1",
x"B4708580",
x"B4D98608",
x"B54C8678",
x"B5C286D2",
x"B639871D",
x"B6B68760",
x"B74087A8",
x"B7E487FB",
x"B8B08862",
x"B9AC88DA",
x"BADC8962",
x"BC3989EF",
x"BDB38A77",
x"BF338AF0",
x"C09D8B4F",
x"C1D78B93",
x"C2CC8BBE",
x"C36E8BDA",
x"C3C38BF7",
x"C3D48C2A",
x"C3BC8C80",
x"C3998D0D",
x"C3898DD5",
x"C3AC8ED9",
x"C412900C",
x"C4C3915B",
x"C5B792AB",
x"C6DE93DF",
x"C81F94DB",
x"C95B9586",
x"CA7795D4",
x"CB5D95BF",
x"CC01954F",
x"CC649497",
x"CC9093AE",
x"CC9892B2",
x"CC9391C2",
x"CC9A90F7",
x"CCBF9063",
x"CD0B9010",
x"CD7F8FFD",
x"CE129022",
x"CEAD906C",
x"CF3D90C7",
x"CFA59118",
x"CFD0914F",
x"CFB39159",
x"CF4A9131",
x"CE9F90D8",
x"CDC79059",
x"CCDB8FC6",
x"CBFC8F38",
x"CB468EC8",
x"CAD08E8B",
x"CAA88E97",
x"CAD08EF4",
x"CB418FA5",
x"CBED90A2",
x"CCBA91DD",
x"CD92933F",
x"CE6094B3",
x"CF13961D",
x"CFA0976B",
x"D0039887",
x"D0409969",
x"D0589A07",
x"D0539A5C",
x"D0369A6B",
x"D0059A33",
x"CFBE99BB",
x"CF629906",
x"CEE89819",
x"CE4A96F9",
x"CD7B95AA",
x"CC6D942E",
x"CB099286",
x"C93690AE",
x"C6D18E9E",
x"C3B48C4F",
x"BFB989B2",
x"BAB986B9",
x"B49E835A",
x"AD607F8E",
x"A5157B5B",
x"9BEC76D0",
x"9235720A",
x"88596D3A",
x"7ED66891",
x"762E6453",
x"6EDC60BB",
x"69455E00",
x"65AD5C49",
x"642D5BAB",
x"64B15C1F",
x"67025D8D",
x"6AC15FC3",
x"6F7D6284",
x"74C2658A",
x"7A216890",
x"7F3E6B5B",
x"83D56DBF",
x"87BF6FA3",
x"8AF370FB",
x"8D7771D1",
x"8F637237",
x"90D37248",
x"91E47223",
x"92AE71DF",
x"933F7195",
x"93A5714F",
x"93E5711A",
x"940070F8",
x"93FB70EC",
x"93DF70F5",
x"93B27113",
x"93817148",
x"93567196",
x"933B71FE",
x"9335727C",
x"9348730F",
x"937173AF",
x"93AE7455",
x"93F674F8",
x"9445758D",
x"9495760C",
x"94E3766F",
x"952B76B6",
x"957076E2",
x"95B376F8",
x"95FA7701",
x"96487705",
x"96A2770D",
x"97147722",
x"97A17747",
x"98547782",
x"993477D2",
x"9A457836",
x"9B8878AA",
x"9CF8792C",
x"9E8E79B6",
x"A0367A44",
x"A1DC7AD6",
x"A3677B64",
x"A4C07BF1",
x"A5D67C78",
x"A69B7CF8",
x"A70D7D71",
x"A7337DDD",
x"A71B7E3A",
x"A6D97E84",
x"A6807EB5",
x"A6267EC7",
x"A5DA7EB9",
x"A5A57E88",
x"A58A7E39",
x"A58A7DD1",
x"A5A27D60",
x"A5D27CF5",
x"A61F7CA9",
x"A68F7C8E",
x"A7327CB9",
x"A8117D3C",
x"A9397E1C",
x"AAB17F57",
x"AC6E80E1",
x"AE63829F",
x"B0718473",
x"B2748638",
x"B43F87C6",
x"B5A88901",
x"B68C89D2",
x"B6DA8A2C",
x"B68A8A14",
x"B5AC8997",
x"B45E88CF",
x"B2C787D7",
x"B11586D0",
x"AF7185D3",
x"ADFF84F3",
x"ACD48439",
x"ABF383A6",
x"AB53832F",
x"AADE82C6",
x"AA7E825E",
x"AA1681ED",
x"A998816A",
x"A8F880DD",
x"A8428050",
x"A7857FD4",
x"A6DE7F82",
x"A66D7F6A",
x"A6497F9B",
x"A6848016",
x"A71F80D4",
x"A80B81C0",
x"A92882BB",
x"AA4783A1",
x"AB38844C",
x"ABCC849F",
x"ABE08485",
x"AB5D83F7",
x"AA4A8300",
x"A8BA81B5",
x"A6D68036",
x"A4CD7EAF",
x"A2D27D3A",
x"A1077BF7",
x"9F847AF1",
x"9E487A25",
x"9D38797E",
x"9C2978DD",
x"9AE4781C",
x"99317718",
x"96DF75B0",
x"93D573D8",
x"90147192",
x"8BB96EF6",
x"87036C2D",
x"823E696B",
x"7DC966E8",
x"7A0064DA",
x"7730636F",
x"759162C1",
x"754462D9",
x"764563B1",
x"787A652D",
x"7BAE6728",
x"7FA0697C",
x"840B6BFC",
x"88AA6E85",
x"8D4370FB",
x"91A97347",
x"95B8755E",
x"995D7737",
x"9C8A78CE",
x"9F3B7A1D",
x"A16B7B20",
x"A31A7BD0",
x"A4437C25",
x"A4E67C1B",
x"A5017BB2",
x"A4977AEF",
x"A3AF79E0",
x"A2567896",
x"A09E7729",
x"9E9E75B4",
x"9C747454",
x"9A3B731C",
x"98117221",
x"9614716E",
x"945D7108",
x"92FE70EB",
x"92097112",
x"91837170",
x"916C71FC",
x"91BE72A7",
x"92697362",
x"93557425",
x"946A74E0",
x"9587758B",
x"9690761F",
x"97697692",
x"97FE76E1",
x"9843770B",
x"9836770D",
x"97DA76EF",
x"973F76B7",
x"9677766E",
x"9594761D",
x"94AC75D1",
x"93CF7592",
x"930A7562",
x"92637548",
x"91DF7543",
x"917E754B",
x"9140755C",
x"9125756F",
x"912E757E",
x"91587581",
x"91A17574",
x"92097557",
x"92837526",
x"930474E5",
x"937D7493",
x"93D77430",
x"940173BD",
x"93E97339",
x"938372A6",
x"92CF7205",
x"91D27158",
x"909F70AA",
x"8F537002",
x"8E0B6F6E",
x"8CEC6EFA",
x"8C146EB8",
x"8B9F6EB4",
x"8B9E6EF5",
x"8C146F7F",
x"8CFA704E",
x"8E3F7155",
x"8FC97282",
x"917973BB",
x"932A74EB",
x"94BB75F5",
x"961276C7",
x"971A7752",
x"97C07792",
x"98047788",
x"97E4773E",
x"976D76C7",
x"96AB7634",
x"95B2759C",
x"949C7510",
x"938074A0",
x"92777455",
x"919D7434",
x"91067440",
x"90C97475",
x"90F174CD",
x"918B7544",
x"929475D4",
x"94077675",
x"95D07722",
x"97D677D4",
x"99F97882",
x"9C127922",
x"9DFE79A8",
x"9F9B7A09",
x"A0CF7A3E",
x"A1877A3E",
x"A1C27A06",
x"A188799D",
x"A0EE790B",
x"A012785D",
x"9F1277A6",
x"9E0D76F7",
x"9D12765D",
x"9C2B75E0",
x"9B4D757E",
x"9A5D752C",
x"993174D4",
x"979A745A",
x"956273A0",
x"925D7289",
x"8E7470FC",
x"89A16EEF",
x"83F96C63",
x"7DB1696F",
x"77146631",
x"708062D9",
x"6A595F9A",
x"65025CA9",
x"60CB5A38",
x"5DEF586B",
x"5C8A5759",
x"5C965702",
x"5DEC575E",
x"604B5850",
x"636659B3",
x"66E65B5C",
x"6A795D22",
x"6DDC5EE3",
x"70DF6081",
x"736C61EF",
x"757F6327",
x"772A642F",
x"788C6514",
x"79CB65E8",
x"7B0A66B5",
x"7C66678E",
x"7DF5687A",
x"7FBB697C",
x"81B86A8F",
x"83DC6BAB",
x"86166CC8",
x"884D6DDB",
x"8A6F6ED8",
x"8C666FBA",
x"8E277079",
x"8FA77117",
x"90E37196",
x"91DC71F8",
x"92937244",
x"930A727B",
x"934672A3",
x"934972BA",
x"931872C1",
x"92B472B4",
x"921E7292",
x"915D7254",
x"907671FC",
x"8F72718A",
x"8E597103",
x"8D3B706C",
x"8C246FCE",
x"8B256F31",
x"8A4C6EA0",
x"89A26E20",
x"892F6DB5",
x"88F46D61",
x"88EF6D20",
x"89156CF0",
x"895D6CCD",
x"89BB6CB1",
x"8A226C9E",
x"8A896C93",
x"8AE76C94",
x"8B3F6CA6",
x"8B906CCF",
x"8BDF6D13",
x"8C346D76",
x"8C946DF3",
x"8D036E85",
x"8D7E6F1E",
x"8E046FB4",
x"8E8B7033",
x"8F07708F",
x"8F6E70BD",
x"8FB770B5",
x"8FD6707A",
x"8FCB7012",
x"8F946F88",
x"8F376EEC",
x"8EBC6E4F",
x"8E2E6DC2",
x"8D976D54",
x"8D006D0C",
x"8C716CEE",
x"8BEF6CF6",
x"8B796D1E",
x"8B0B6D5E",
x"8AA46DA4",
x"8A3C6DE6",
x"89CF6E17",
x"89566E30",
x"88D06E29",
x"883F6E00",
x"87A56DBB",
x"87066D5C",
x"86696CEC",
x"85D66C73",
x"854F6BF8",
x"84D96B7C",
x"84736B04",
x"84156A8D",
x"83BB6A14",
x"83586993",
x"82E26904",
x"82536866",
x"81A567BA",
x"80D96701",
x"7FF76649",
x"7F0A65A0",
x"7E246511",
x"7D5564AF",
x"7CAE6486",
x"7C39649B",
x"7BFD64F2",
x"7BF4657D",
x"7C166631",
x"7C4F66F5",
x"7C8B67AE",
x"7CB56845",
x"7CB568A3",
x"7C7F68B5",
x"7C076875",
x"7B4B67E0",
x"7A4C6700",
x"791065E3",
x"77A06498",
x"76016335",
x"743D61C6",
x"72516058",
x"70445EF3",
x"6E195D98",
x"6BD55C48",
x"69825B02",
x"672E59C6",
x"64F05895",
x"62E15777",
x"611A5677",
x"5FB455A1",
x"5EC55505",
x"5E5B54B0",
x"5E7954AD",
x"5F1C5505",
x"603455B6",
x"61AD56BC",
x"636D580A",
x"655C5991",
x"67645B40",
x"69705D04",
x"6B765ECD",
x"6D706088",
x"6F5C6229",
x"713C63A4",
x"731764F3",
x"74F0660E",
x"76CC66F6",
x"78AB67AB",
x"7A8D6831",
x"7C6D688D",
x"7E4468CB",
x"800968F3",
x"81B26913",
x"83356934",
x"848A6962",
x"85A769A0",
x"868769F3",
x"872C6A5B",
x"879B6AD2",
x"87DB6B54",
x"87FA6BD7",
x"880A6C54",
x"881A6CC8",
x"88396D2D",
x"88766D85",
x"88D26DCD",
x"894E6E08",
x"89D96E37",
x"8A666E58",
x"8ADA6E68",
x"8B1D6E62",
x"8B176E43",
x"8AB86E00",
x"89F76D9A",
x"88D96D0F",
x"876D6C61",
x"85CB6B99",
x"84146AC4",
x"826C69EF",
x"80F4692A",
x"7FCC6883",
x"7F0A6807",
x"7EBA67BE",
x"7ED967AA",
x"7F6067C9",
x"80386817",
x"8148688C",
x"826F691B",
x"838D69BB",
x"84876A5E",
x"85456AF9",
x"85B46B80",
x"85CF6BE8",
x"85946C28",
x"850E6C37",
x"844F6C10",
x"836C6BB2",
x"82806B24",
x"81A86A6D",
x"80FE69A0",
x"809668D1",
x"807E6816",
x"80BF678A",
x"81556741",
x"82376749",
x"835267AA",
x"8491685F",
x"85DC6959",
x"871A6A83",
x"88376BBE",
x"89216CEE",
x"89CF6DF3",
x"8A3B6EBA",
x"8A676F34",
x"8A5A6F5F",
x"8A1B6F43",
x"89B56EEE",
x"89346E75",
x"889F6DF0",
x"88066D75",
x"876C6D13",
x"86DB6CD1",
x"86596CB1",
x"85ED6CAB",
x"859E6CB5",
x"856F6CBE",
x"855C6CBA",
x"85656C9C",
x"85836C5E",
x"85AA6C00",
x"85CC6B87",
x"85DB6B00",
x"85C66A75",
x"858169F0",
x"85036980",
x"84496928",
x"835868EB",
x"823968C7",
x"810068B4",
x"7FBF68AA",
x"7E8B689E",
x"7D796889",
x"7C976863",
x"7BEC682A",
x"7B7A67DB",
x"7B37677A",
x"7B0E670A",
x"7AEC668E",
x"7AB2660D",
x"7A446584",
x"798A64F4",
x"7870645C",
x"76F063B8",
x"750D6304",
x"72D8623E",
x"706C6169",
x"6DEE6086",
x"6B865F9B",
x"69615EB3",
x"67A45DD7",
x"666C5D14",
x"65CB5C73",
x"65C75BFA",
x"66565BB3",
x"67685BA1",
x"68E15BC3",
x"6AA15C1C",
x"6C905CA9",
x"6E965D6A",
x"70A35E5C",
x"72B15F7D",
x"74C260CC",
x"76DF6241",
x"790E63D6",
x"7B5B6583",
x"7DC86737",
x"805868E5",
x"82FE6A7C",
x"85B26BEC",
x"885C6D27",
x"8AEA6E24",
x"8D456EDE",
x"8F596F54",
x"911A6F90",
x"927E6F9F",
x"93876F8F",
x"943C6F76",
x"94AC6F68",
x"94EC6F76",
x"95156FAE",
x"9545701C",
x"959070C0",
x"960A7195",
x"96BC728F",
x"97A2739C",
x"98A974A0",
x"99AF7581",
x"9A85761F",
x"9AF47660",
x"9AC5762A",
x"99C37572",
x"97CF7433",
x"94D77275",
x"90EC704E",
x"8C346DD9",
x"86F06B3F",
x"817368AA",
x"7C1B6641",
x"77426428",
x"7338627C",
x"70376149",
x"6E586097",
x"6D9E6059",
x"6DEA607D",
x"6F0A60EA",
x"70BC6183",
x"72B86228",
x"74BB62C1",
x"768B633B",
x"7800638A",
x"790163A8",
x"798A6398",
x"79A46365",
x"7960631A",
x"78DB62C8",
x"782D6280",
x"7770624F",
x"76BA623F",
x"76136258",
x"75836297",
x"750A62F4",
x"749E6365",
x"743463D3",
x"73BF642A",
x"73326455",
x"7287643F",
x"71BE63E0",
x"70DC6334",
x"6FF66246",
x"6F28612D",
x"6E996008",
x"6E705F06",
x"6ED95E4F",
x"6FF65E10",
x"71DB5E67",
x"748E5F69",
x"78016115",
x"7C10635C",
x"80836617",
x"85186914",
x"89846C1C",
x"8D806EEF",
x"90CE715A",
x"93437333",
x"94C97461",
x"956474E0",
x"952C74BB",
x"94507415",
x"93057313",
x"918A71E4",
x"901870B4",
x"8EDF6FA7",
x"8DFD6ED8",
x"8D836E54",
x"8D6D6E17",
x"8DAA6E19",
x"8E1E6E44",
x"8EA86E82",
x"8F2B6EBE",
x"8F8E6EE9",
x"8FBF6EFA",
x"8FB96EF0",
x"8F816ED1",
x"8F246EA7",
x"8EAE6E80",
x"8E2E6E66",
x"8DAC6E5E",
x"8D286E65",
x"8C9A6E6E",
x"8BEC6E68",
x"8B036E38",
x"89BE6DC2",
x"87FE6CEC",
x"85AC6BA1",
x"82B769D5",
x"7F1E6787",
x"7AF364C6",
x"765561AE",
x"71725E64",
x"6C805B1A",
x"67BF57FE",
x"63695542",
x"5FB3530B",
x"5CC75178",
x"5AC25096",
x"59B05068",
x"598950DE",
x"5A3D51DD",
x"5BAA5343",
x"5DA954ED",
x"600D56B3",
x"62A8587A",
x"65515A25",
x"67DF5BA8",
x"6A355CF7",
x"6C3E5E12",
x"6DEC5EFD",
x"6F3B5FBB",
x"70316050",
x"70D960C5",
x"7147611B",
x"718E6156",
x"71C86179",
x"720A6188",
x"7266618B",
x"72E96184",
x"7397617D",
x"746D6176",
x"75606173",
x"765C6172",
x"774C616D",
x"7816615C",
x"78A46135",
x"78E560F2",
x"78CF608A",
x"78606000",
x"77A35F59",
x"76A45EA5",
x"757D5DF3",
x"74495D59",
x"73215CE9",
x"721E5CB2",
x"71525CBD",
x"70CB5D0B",
x"708C5D91",
x"70915E41",
x"70D15F06",
x"713C5FCB",
x"71C2607E",
x"72536110",
x"72E06176",
x"735E61B2",
x"73C561C6",
x"741461BE",
x"744E61A1",
x"7474617D",
x"74906159",
x"74A3613B",
x"74B26124",
x"74BE6113",
x"74C56104",
x"74C260F4",
x"74B260E2",
x"748E60CB",
x"745560B4",
x"740760A1",
x"73AB609B",
x"734B60AB",
x"72F360D5",
x"72B4611D",
x"729D6181",
x"72BD61FE",
x"7317628B",
x"73AD631A",
x"7474639A",
x"755E63FD",
x"76506437",
x"7735643C",
x"77F2640E",
x"787063AD",
x"78A76321",
x"7894627A",
x"784261CC",
x"77C46128",
x"773860A4",
x"76BC604F",
x"76736035",
x"7673605C",
x"76D160C5",
x"778D6168",
x"78A26238",
x"79FD6327",
x"7B7F6425",
x"7D076521",
x"7E75660A",
x"7FA866D5",
x"808D6779",
x"811A67F2",
x"814C683B",
x"81316859",
x"80D9684E",
x"805B681E",
x"7FCC67D2",
x"7F44676D",
x"7ED266F9",
x"7E7D667A",
x"7E4B65FA",
x"7E32657F",
x"7E2E650E",
x"7E3064AF",
x"7E2A6468",
x"7E13643B",
x"7DDF642B",
x"7D8A6435",
x"7D116458",
x"7C74648B",
x"7BB564C6",
x"7AD264FD",
x"79CF6524",
x"78A8652D",
x"775C650A",
x"75E964B5",
x"74496427",
x"7280635C",
x"70916259",
x"6E866128",
x"6C6F5FD8",
x"6A635E78",
x"687C5D24",
x"66D95BEE",
x"65965AEE",
x"64CD5A35",
x"649059D2",
x"64E659C9",
x"65D15A1B",
x"673E5AC2",
x"69195BAC",
x"6B3F5CC8",
x"6D935E00",
x"6FEF5F3B",
x"72356067",
x"744F6173",
x"762D6253",
x"77CB6301",
x"792A6380",
x"7A5563D6",
x"7B596411",
x"7C46643E",
x"7D2A6470",
x"7E0E64B7",
x"7EFC651E",
x"7FF365B2",
x"80F76677",
x"8201676C",
x"83106889",
x"841D69C1",
x"85216B04",
x"861B6C41",
x"87036D65",
x"87D66E5C",
x"88906F1E",
x"89296FA0",
x"899E6FDF",
x"89E76FDE",
x"89FE6FA6",
x"89E06F41",
x"898B6EBA",
x"89016E1E",
x"88486D79",
x"87696CD5",
x"86716C38",
x"85716BA7",
x"847A6B24",
x"839E6AB4",
x"82ED6A55",
x"82746A0A",
x"823B69D4",
x"824669B2",
x"829369A6",
x"831B69B0",
x"83D369CF",
x"84AE6A06",
x"859A6A4F",
x"86886AAD",
x"87696B1C",
x"88346B9A",
x"88DF6C24",
x"89696CB7",
x"89D26D4E",
x"8A1D6DE1",
x"8A506E6B",
x"8A746EE1",
x"8A8D6F3E",
x"8AA16F7A",
x"8AB56F92",
x"8AC96F83",
x"8ADF6F4F",
x"8AF36EFA",
x"8B036E90",
x"8B076E16",
x"8AFD6D99",
x"8AE06D23",
x"8AAE6CBA",
x"8A636C63",
x"8A036C23",
x"898D6BF5",
x"890B6BDB",
x"88836BCC",
x"87FD6BCA",
x"87846BCE",
x"87226BDB",
x"86DC6BED",
x"86B86C0C",
x"86B56C37",
x"86D56C75",
x"870E6CC8",
x"875D6D31",
x"87B86DB1",
x"88186E45",
x"88776EE6",
x"88D36F8F",
x"892B7035",
x"898470D1",
x"89E37158",
x"8A4C71C3",
x"8AC6720C",
x"8B537230",
x"8BF47231",
x"8CA57210",
x"8D5F71D4",
x"8E187186",
x"8EC97131",
x"8F6470DF",
x"8FE4709A",
x"90437069",
x"907C7051",
x"908E7052",
x"907C706B",
x"90497093",
x"8FF970C4",
x"8F9070EF",
x"8F10710A",
x"8E7A710C",
x"8DCF70EC",
x"8D0A70A3",
x"8C27702E",
x"8B1A6F8C",
x"89DA6EBA",
x"88586DB7",
x"86846C83",
x"844E6B19",
x"81AA6976",
x"7E8E679A",
x"7AFD6583",
x"7704633B",
x"72BB60CE",
x"6E4C5E4F",
x"69E95BDD",
x"65CE599A",
x"623B57A6",
x"5F695623",
x"5D8C552E",
x"5CC054D0",
x"5D105512",
x"5E7055E7",
x"60BB5738",
x"63BD58E6",
x"67345ACA",
x"6ADB5CC3",
x"6E735EAF",
x"71C76076",
x"74B2620A",
x"77246366",
x"791B648B",
x"7AA56583",
x"7BDE6656",
x"7CDF670E",
x"7DC567B1",
x"7EA8683F",
x"7F9768BB",
x"809D6924",
x"81BC6979",
x"82F669BE",
x"844969FC",
x"85B66A3B",
x"87436A8D",
x"88F26AFF",
x"8AC86BA0",
x"8CCC6C78",
x"8EFC6D89",
x"91536ED1",
x"93C67044",
x"964371D5",
x"98B47371",
x"9B007503",
x"9D11767C",
x"9ED377CE",
x"A03B78EE",
x"A14379D8",
x"A1EE7A8C",
x"A2467B0B",
x"A25C7B57",
x"A23F7B77",
x"A2047B71",
x"A1BB7B4A",
x"A1737B0C",
x"A13B7AC0",
x"A11B7A6F",
x"A11B7A28",
x"A14379F5",
x"A19B79E7",
x"A2257A08",
x"A2E77A5D",
x"A3E47AEB",
x"A5197BAC",
x"A6807C98",
x"A8077D9B",
x"A99E7EA0",
x"AB287F92",
x"AC8A8059",
x"ADA880E1",
x"AE6A811E",
x"AEC2810A",
x"AEAC80A9",
x"AE308008",
x"AD677F3F",
x"AC707E65",
x"AB6D7D96",
x"AA877CEA",
x"A9DF7C75",
x"A9887C43",
x"A98A7C56",
x"A9D97CA2",
x"AA5D7D18",
x"AAF37DA3",
x"AB6B7E28",
x"ABA17E8F",
x"AB6E7EC6",
x"AABF7EBF",
x"A9877E75",
x"A7D07DED",
x"A5B17D2D",
x"A34B7C49",
x"A0C37B4E",
x"9E467A51",
x"9BF7795D",
x"99F7787F",
x"985A77BC",
x"97317716",
x"967D768F",
x"963C7625",
x"966475D4",
x"96E4759C",
x"97A9757B",
x"989A7571",
x"999C757E",
x"9A94759F",
x"9B6475D0",
x"9BF7760F",
x"9C337651",
x"9C10768D",
x"9B8376BC",
x"9A9276CE",
x"994C76C0",
x"97C27688",
x"96117623",
x"94537595",
x"92A274E0",
x"9115740C",
x"8FBF7326",
x"8EA7723B",
x"8DD2715B",
x"8D3C7094",
x"8CDF6FF5",
x"8CAC6F86",
x"8C956F4F",
x"8C8A6F51",
x"8C796F85",
x"8C4E6FDC",
x"8BF47045",
x"8B5870A4",
x"8A6670DE",
x"891070D2",
x"8749706B",
x"850E6F94",
x"82666E45",
x"7F5F6C83",
x"7C116A5B",
x"78A167EB",
x"75376556",
x"720062C8",
x"6F2A606A",
x"6CE05E67",
x"6B445CE0",
x"6A725BED",
x"6A765B9B",
x"6B575BED",
x"6D0C5CD9",
x"6F865E50",
x"72AD603C",
x"76656286",
x"7A8E6510",
x"7F0D67C2",
x"83C26A86",
x"88906D45",
x"8D5D6FEB",
x"92117266",
x"969574AA",
x"9AD276AC",
x"9EB17861",
x"A21E79C6",
x"A5077AD8",
x"A75C7B9B",
x"A9147C12",
x"AA2B7C44",
x"AAA17C3D",
x"AA807C05",
x"A9DA7BA5",
x"A8C97B26",
x"A7647A92",
x"A5CF79F1",
x"A428794A",
x"A28E78A7",
x"A11F7816",
x"9FF477A0",
x"9F227757",
x"9EBC7744",
x"9ECF7774",
x"9F6377EF",
x"A07A78B7",
x"A21479C7",
x"A4247B16",
x"A69B7C92",
x"A9637E26",
x"AC5E7FBC",
x"AF6B8140",
x"B26D82A2",
x"B54283D9",
x"B7D184E0",
x"BA0885BF",
x"BBE08681",
x"BD598736",
x"BE7887F1",
x"BF4D88BB",
x"BFE3899B",
x"C0448A90",
x"C0778B8A",
x"C07B8C79",
x"C04D8D42",
x"BFE38DCC",
x"BF398E04",
x"BE4C8DDC",
x"BD268D53",
x"BBDD8C76",
x"BA8F8B5A",
x"B9678A27",
x"B89288FE",
x"B83A8808",
x"B8828767",
x"B978872F",
x"BB1C8767",
x"BD50880B",
x"BFEA8904",
x"C2AD8A35",
x"C5598B7B",
x"C7AB8CB2",
x"C96F8DB9",
x"CA7F8E79",
x"CACD8EE3",
x"CA5D8EF6",
x"C94A8EB7",
x"C7BA8E35",
x"C5DE8D86",
x"C3EA8CBE",
x"C2098BF4",
x"C0648B3F",
x"BF128AAE",
x"BE238A4D",
x"BD998A27",
x"BD6F8A39",
x"BD988A84",
x"BE018AFD",
x"BE958B98",
x"BF418C43",
x"BFEE8CED",
x"C08B8D81",
x"C1078DF1",
x"C1568E32",
x"C1708E3C",
x"C1578E14",
x"C10F8DC1",
x"C0A18D4C",
x"C0188CC6",
x"BF7F8C3C",
x"BEE08BB6",
x"BE398B3B",
x"BD858AC8",
x"BCBA8A56",
x"BBC389DC",
x"BA8E8950",
x"B90B88A9",
x"B72D87E9",
x"B4F8870D",
x"B2758621",
x"AFBC8531",
x"ACE78443",
x"AA128361",
x"A754828A",
x"A4BB81B0",
x"A23F80C0",
x"9FCF7FA0",
x"9D427E33",
x"9A6D7C59",
x"971D79FF",
x"932A771F",
x"8E7A73C3",
x"890E7003",
x"82FE6C06",
x"7C8167FD",
x"75E2641E",
x"6F79609B",
x"69A75D9C",
x"64BF5B40",
x"610A5991",
x"5EB1588F",
x"5DC0582B",
x"5E245847",
x"5FB158CA",
x"62285994",
x"653B5A87",
x"689A5B8B",
x"6BFF5C91",
x"6F2E5D8B",
x"71FF5E77",
x"745E5F4F",
x"76466017",
x"77C660CE",
x"78F6617A",
x"79EC621D",
x"7AC762BC",
x"7B9A635F",
x"7C766407",
x"7D5E64BA",
x"7E4F657A",
x"7F416648",
x"8027671E",
x"80F267F7",
x"819668C8",
x"820B6984",
x"82506A23",
x"826C6A9A",
x"82666AE6",
x"824C6B07",
x"822F6B03",
x"821E6AE3",
x"82246AB7",
x"82486A89",
x"828B6A68",
x"82EC6A5B",
x"83606A68",
x"83DD6A8C",
x"845C6AC1",
x"84D06B00",
x"85366B3E",
x"858D6B72",
x"85D96B90",
x"86216B96",
x"866C6B80",
x"86C36B4F",
x"87316B0A",
x"87B56AB8",
x"88556A62",
x"890B6A10",
x"89D669CF",
x"8AAB69A8",
x"8B8369A3",
x"8C5369C4",
x"8D116A10",
x"8DB46A87",
x"8E346B26",
x"8E8B6BE5",
x"8EB86CBE",
x"8EB76DA6",
x"8E8D6E90",
x"8E416F73",
x"8DDD7047",
x"8D707103",
x"8D0771A4",
x"8CB47229",
x"8C837290",
x"8C7B72DB",
x"8CA5730D",
x"8CF97326",
x"8D6F7329",
x"8DF47316",
x"8E7972EC",
x"8EE472AD",
x"8F29725B",
x"8F3871F9",
x"8F0D718C",
x"8EAB711A",
x"8E1E70AB",
x"8D797048",
x"8CD26FF8",
x"8C3C6FBD",
x"8BCF6F9A",
x"8B936F8D",
x"8B8D6F92",
x"8BB56F9F",
x"8C006FA9",
x"8C566FA7",
x"8CA16F92",
x"8CCC6F62",
x"8CC66F16",
x"8C846EB0",
x"8C0A6E37",
x"8B5F6DB5",
x"8A976D38",
x"89CE6CCE",
x"891D6C7F",
x"889F6C54",
x"886A6C51",
x"888A6C76",
x"88FD6CBD",
x"89BC6D1D",
x"8AB46D8C",
x"8BC86E00",
x"8CD96E72",
x"8DC86ED9",
x"8E7C6F34",
x"8EDC6F85",
x"8EE06FCD",
x"8E847010",
x"8DD27054",
x"8CD87096",
x"8BA770D5",
x"8A56710C",
x"88F3712D",
x"8788712B",
x"861770F5",
x"84977078",
x"82F36FA6",
x"81176E72",
x"7EE76CD8",
x"7C4F6AD7",
x"79426879",
x"75BE65D0",
x"71D562F6",
x"6DA5600D",
x"695F5D35",
x"653B5A97",
x"61785854",
x"5E4F568C",
x"5BF55554",
x"5A8D54B9",
x"5A2754BA",
x"5AC0554D",
x"5C41565E",
x"5E8457D0",
x"61595981",
x"648C5B52",
x"67E65D1F",
x"6B3B5ED3",
x"6E66605C",
x"715161AE",
x"73EC62CC",
x"763563B9",
x"78346486",
x"79F2653F",
x"7B8065F3",
x"7CED66B1",
x"7E496781",
x"7FA46869",
x"81046966",
x"82736A72",
x"83EF6B83",
x"85746C8A",
x"86FD6D7C",
x"887A6E4A",
x"89DD6EE6",
x"8B156F4E",
x"8C146F7A",
x"8CCF6F6F",
x"8D416F31",
x"8D676ECB",
x"8D4F6E48",
x"8D046DBA",
x"8C9A6D2D",
x"8C246CB0",
x"8BB66C51",
x"8B626C16",
x"8B346C0A",
x"8B316C2E",
x"8B596C83",
x"8BAA6D08",
x"8C1E6DB5",
x"8CAF6E85",
x"8D5C6F6B",
x"8E20705F",
x"8F007154",
x"9001723E",
x"91287316",
x"927A73D5",
x"93F97478",
x"959F74FF",
x"9767756E",
x"994075CB",
x"9B15761F",
x"9CD2766E",
x"9E5C76C0",
x"9F9F7718",
x"A08B7771",
x"A11877C8",
x"A1457819",
x"A118785A",
x"A0A27882",
x"9FF7788F",
x"9F327881",
x"9E6E785B",
x"9DC87825",
x"9D5277EC",
x"9D1E77BD",
x"9D3577A3",
x"9D9577A7",
x"9E3577CB",
x"9F03780D",
x"9FEA7868",
x"A0D078CD",
x"A19C7932",
x"A23C7986",
x"A29E79C3",
x"A2BC79E0",
x"A29879DD",
x"A23D79C0",
x"A1BC7990",
x"A12B795A",
x"A0A17928",
x"A02E7902",
x"9FE378EF",
x"9FC678EF",
x"9FD078FC",
x"9FF4790B",
x"A01F790F",
x"A03578FC",
x"A01B78C3",
x"9FBC785B",
x"9F0777C4",
x"9DF876FF",
x"9C9B761C",
x"9B037527",
x"994F743B",
x"97A8736E",
x"963872D4",
x"9524727E",
x"94867275",
x"946C72B6",
x"94D37337",
x"95A473E6",
x"96BD74AA",
x"97F17567",
x"990E7602",
x"99E97667",
x"9A5F768B",
x"9A59766A",
x"99D6760B",
x"98E2757B",
x"979874CB",
x"9617740D",
x"947E7350",
x"92EA7297",
x"916471E1",
x"8FED7124",
x"8E74704F",
x"8CDF6F51",
x"8B0B6E14",
x"88DD6C92",
x"86436AC7",
x"833968BC",
x"7FD26687",
x"7C2F6446",
x"7889621B",
x"751A602B",
x"72245E95",
x"6FDF5D74",
x"6E765CD7",
x"6DFF5CC3",
x"6E785D36",
x"6FCC5E1F",
x"71D35F6D",
x"745C610A",
x"772E62DF",
x"7A1464D5",
x"7CE666D9",
x"7F8468DB",
x"81E06ACB",
x"83FA6C9D",
x"85DC6E47",
x"87976FBD",
x"893F70FC",
x"8AE97200",
x"8CA172CB",
x"8E6C735F",
x"904573C6",
x"92217408",
x"93F07431",
x"959B7451",
x"9710746F",
x"983E7493",
x"991F74C6",
x"99B27506",
x"9A047558",
x"9A2475B7",
x"9A297622",
x"9A2F7699",
x"9A4D771B",
x"9A9A77A6",
x"9B1E783D",
x"9BDD78DD",
x"9CD67985",
x"9DF87A30",
x"9F387AD8",
x"A0807B79",
x"A1C87C0E",
x"A3057C94",
x"A43B7D08",
x"A5747D74",
x"A6BF7DDD",
x"A82E7E4D",
x"A9D17ED0",
x"ABB57F6D",
x"ADDA802D",
x"B039810F",
x"B2BC820C",
x"B547831C",
x"B7B6842D",
x"B9E68533",
x"BBB6861C",
x"BD1286DE",
x"BDEE8771",
x"BE4C87D4",
x"BE378808",
x"BDC98818",
x"BD1F880B",
x"BC5687EE",
x"BB8F87CD",
x"BAE487B3",
x"BA6A87AB",
x"BA3287BB",
x"BA4487EC",
x"BAA88842",
x"BB6088C2",
x"BC6A896F",
x"BDC38A43",
x"BF658B3E",
x"C1498C52",
x"C35E8D74",
x"C5958E97",
x"C7D68FAA",
x"CA0790A0",
x"CC0E916D",
x"CDD09210",
x"CF319283",
x"D01F92CE",
x"D08B92F4",
x"D06B9302",
x"CFC392F9",
x"CE9C92E0",
x"CD0892B9",
x"CB1E927D",
x"C8F89228",
x"C6B591B2",
x"C4719114",
x"C244904C",
x"C0478F5C",
x"BE858E4C",
x"BD058D27",
x"BBC98BFE",
x"BACA8AE4",
x"B9FF89EC",
x"B9608922",
x"B8DE8891",
x"B872883F",
x"B8148829",
x"B7C08848",
x"B772888D",
x"B72B88E7",
x"B6E48943",
x"B69E898E",
x"B65189B4",
x"B5FD89A7",
x"B59B895F",
x"B52E88DA",
x"B4B98821",
x"B44A8740",
x"B3EE8650",
x"B3B58566",
x"B3AC849B",
x"B3D98401",
x"B430839F",
x"B4998370",
x"B4E8835D",
x"B4E18345",
x"B43C82F7",
x"B2B58242",
x"B00C80F4",
x"AC1F7EED",
x"A6DE7C15",
x"A0667877",
x"98F37430",
x"90E36F79",
x"88AA6A99",
x"80C365E2",
x"79A861A7",
x"73BB5E2E",
x"6F445BAB",
x"6C635A38",
x"6B1959D6",
x"6B3D5A6B",
x"6C945BCC",
x"6ED15DBF",
x"71A3600A",
x"74C16274",
x"77F064D0",
x"7B096701",
x"7DF668F7",
x"80B56AB0",
x"83506C34",
x"85D86D92",
x"885C6ED4",
x"8AE77006",
x"8D80712D",
x"901F7245",
x"92BE7348",
x"9546742F",
x"97A874EC",
x"99D3757E",
x"9BBE75E4",
x"9D647623",
x"9ECD764B",
x"A004766C",
x"A11C769B",
x"A22976E5",
x"A33F775D",
x"A46E7809",
x"A5BC78ED",
x"A72B7A03",
x"A8B07B43",
x"AA3D7C9B",
x"ABBF7DFC",
x"AD1C7F54",
x"AE468095",
x"AF2B81AD",
x"AFC28295",
x"B00C8342",
x"B01283B3",
x"AFE083EA",
x"AF8883EA",
x"AF1F83BB",
x"AEB68367",
x"AE6082FD",
x"AE26828B",
x"AE128221",
x"AE2881CD",
x"AE64819F",
x"AEC681A2",
x"AF4A81DC",
x"AFEB824C",
x"B0A582F0",
x"B17283BD",
x"B25084A3",
x"B33A8592",
x"B42D8673",
x"B5238732",
x"B61887BF",
x"B707880E",
x"B7EB881D",
x"B8C187EC",
x"B987878A",
x"BA3A8708",
x"BADD8680",
x"BB71860A",
x"BBFB85C2",
x"BC8485BB",
x"BD128605",
x"BDB086A7",
x"BE67879B",
x"BF3C88D6",
x"C0358A43",
x"C1508BC9",
x"C2888D4E",
x"C3D38EB8",
x"C5238FF3",
x"C66790F3",
x"C78C91B1",
x"C881922E",
x"C9399270",
x"C9A99282",
x"C9CA926C",
x"C99B9238",
x"C91F91E9",
x"C85A9182",
x"C75190FD",
x"C60C9055",
x"C48F8F84",
x"C2E18E87",
x"C1078D5C",
x"BF0C8C08",
x"BCFE8A9D",
x"BAED8925",
x"B8F187BC",
x"B7268678",
x"B5A5856E",
x"B48584B2",
x"B3DA844A",
x"B3AB8438",
x"B3F08474",
x"B49884EC",
x"B57F8584",
x"B67F8622",
x"B76886A8",
x"B80E86FE",
x"B8478711",
x"B7FE86D6",
x"B725864D",
x"B5C28580",
x"B3E7847A",
x"B1B38350",
x"AF468216",
x"ACBD80D9",
x"AA2F7FA0",
x"A7A57E6D",
x"A5197D33",
x"A27D7BE4",
x"9FB37A6D",
x"9CA478B9",
x"993476BA",
x"9556746C",
x"910E71D8",
x"8C736F0F",
x"87A86C2E",
x"82E4695F",
x"7E6766CB",
x"7A6D6497",
x"772B62E4",
x"74C861C6",
x"7356613F",
x"72D26146",
x"732461C5",
x"74206298",
x"7594639E",
x"774664AF",
x"790665B1",
x"7AAB6690",
x"7C1D6744",
x"7D5267CF",
x"7E566844",
x"7F3C68B2",
x"80226930",
x"812769CF",
x"82656A9C",
x"83ED6B99",
x"85CB6CC1",
x"87F96E06",
x"8A6C6F59",
x"8D1070A3",
x"8FCC71D4",
x"928872DE",
x"952E73BA",
x"97AC7468",
x"99F774EE",
x"9C08755A",
x"9DDF75B9",
x"9F7A7617",
x"A0DD7683",
x"A20D7703",
x"A30E779B",
x"A3E77848",
x"A4A17905",
x"A54379CA",
x"A5DC7A8F",
x"A67A7B4D",
x"A7297BFF",
x"A7FA7CA2",
x"A8F77D36",
x"AA2B7DBD",
x"AB987E3D",
x"AD3F7EB9",
x"AF1F7F35",
x"B1307FB6",
x"B36D803F",
x"B5CA80D1",
x"B846816B",
x"BAD7820F",
x"BD7D82BB",
x"C02D836B",
x"C2E18423",
x"C58B84E1",
x"C81C85A3",
x"CA81866C",
x"CCA08736",
x"CE678805",
x"CFC188D9",
x"D0A389AF",
x"D10B8A85",
x"D0F98B59",
x"D07E8C2A",
x"CFAC8CEF",
x"CE988DA7",
x"CD5E8E49",
x"CC108ECF",
x"CAC38F31",
x"C97E8F67",
x"C8478F6C",
x"C71D8F38",
x"C5FC8EC9",
x"C4DB8E1D",
x"C3B68D36",
x"C2888C1D",
x"C1548AD9",
x"C01F897B",
x"BEF78815",
x"BDED86B9",
x"BD148580",
x"BC7E847D",
x"BC4083C0",
x"BC638357",
x"BCE88349",
x"BDC7838F",
x"BEE88421",
x"C02C84E4",
x"C16485BF",
x"C260868E",
x"C2EF8731",
x"C2EB8788",
x"C239877D",
x"C0D18707",
x"BEC18627",
x"BC3084EE",
x"B953837B",
x"B66B81F1",
x"B3C0807B",
x"B1917F40",
x"B00F7E64",
x"AF567DF8",
x"AF697E04",
x"B02E7E7F",
x"B17B7F51",
x"B314805B",
x"B4B28171",
x"B615826A",
x"B708831E",
x"B7658371",
x"B71C8352",
x"B63582BC",
x"B4C681BC",
x"B2F58068",
x"B0F17EE0",
x"AEE67D41",
x"ACF47BB0",
x"AB337A47",
x"A9A67918",
x"A8437829",
x"A6EE7774",
x"A58276E8",
x"A3DA7671",
x"A1D275EF",
x"9F53754B",
x"9C55746E",
x"98E4734A",
x"951E71DE",
x"912E7034",
x"8D4D6E63",
x"89B56C84",
x"869A6ABB",
x"84256927",
x"827067E5",
x"817E6709",
x"814366A0",
x"81A566AA",
x"827A671E",
x"839D67ED",
x"84E36900",
x"86316A3F",
x"87736B96",
x"88A16CEF",
x"89BF6E3D",
x"8ADA6F78",
x"8C03709C",
x"8D4D71AB",
x"8EC872AF",
x"907E73AC",
x"927974AC",
x"94B975B9",
x"973F76D8",
x"9A077810",
x"9D0E7964",
x"A04A7AD6",
x"A3B67C61",
x"A7457E04",
x"AAE37FB5",
x"AE7A8172",
x"B1F28331",
x"B52B84E4",
x"B8018685",
x"BA578804",
x"BC158956",
x"BD298A6D",
x"BD8F8B3C",
x"BD508BB8",
x"BC828BD8",
x"BB468B98",
x"B9C28AFA",
x"B8238A04",
x"B69588C9",
x"B53D8760",
x"B43D85E7",
x"B3AB8481",
x"B38F8352",
x"B3F38278",
x"B4CA8211",
x"B6098226",
x"B7A082BD",
x"B97783CA",
x"BB758532",
x"BD8486D4",
x"BF898888",
x"C1728A22",
x"C3298B80",
x"C49F8C83",
x"C5C98D1D",
x"C6A28D49",
x"C7278D14",
x"C7618C93",
x"C7578BE2",
x"C71C8B1D",
x"C6BD8A62",
x"C64E89C3",
x"C5E3894D",
x"C5858903",
x"C54388DA",
x"C51F88C6",
x"C51B88B4",
x"C52D8894",
x"C54D8859",
x"C56E87FB",
x"C5818781",
x"C57B86F1",
x"C551865C",
x"C50285D4",
x"C48C856D",
x"C3F98535",
x"C3518533",
x"C2A6856C",
x"C20485D4",
x"C1788660",
x"C10E86FB",
x"C0C68791",
x"C09D880E",
x"C08C8862",
x"C07E8884",
x"C0638871",
x"C020882F",
x"BFA387C6",
x"BEDB873F",
x"BDBC86A9",
x"BC42860E",
x"BA748574",
x"B85E84E3",
x"B619845A",
x"B3BF83D9",
x"B1708360",
x"AF4782ED",
x"AD638281",
x"ABD9821E",
x"AAB381C5",
x"A9F68178",
x"A99A8139",
x"A98B8102",
x"A9B280D1",
x"A9F1809C",
x"AA28805B",
x"AA3C8005",
x"AA157F94",
x"A9A97F02",
x"A8F77E59",
x"A8057D98",
x"A6E47CCC",
x"A5A77BFF",
x"A45F7B39",
x"A3187A7C",
x"A1D079C3",
x"A07A7901",
x"9EFD7820",
x"9D327709",
x"9AF175A3",
x"981173D8",
x"9474719C",
x"900B6EEE",
x"8ADF6BDC",
x"850B6881",
x"7EC66504",
x"78586194",
x"72115E62",
x"6C485B9B",
x"67485963",
x"634E57D4",
x"608256F8",
x"5EEC56C9",
x"5E825733",
x"5F1C5818",
x"60805953",
x"62725AB9",
x"64AD5C26",
x"66F55D76",
x"691D5E8D",
x"6B065F5F",
x"6CA65FE3",
x"6DFD6022",
x"6F236027",
x"702E6007",
x"713E5FDA",
x"726C5FBE",
x"73CC5FC6",
x"75666007",
x"773A608B",
x"79386159",
x"7B4E6269",
x"7D5F63B1",
x"7F4F651B",
x"81086694",
x"82766801",
x"838B694E",
x"84496A66",
x"84B56B3D",
x"84DD6BCC",
x"84D26C16",
x"84AA6C20",
x"84776BF9",
x"84496BB0",
x"842B6B57",
x"84226AFC",
x"842E6AAD",
x"84486A72",
x"84696A4C",
x"84896A38",
x"849D6A30",
x"84A26A2A",
x"84956A1D",
x"847C6A06",
x"845C69E1",
x"844469B5",
x"84426990",
x"84666980",
x"84BF6999",
x"855B69EB",
x"863B6A84",
x"87636B69",
x"88C86C96",
x"8A586DF6",
x"8BFE6F73",
x"8D9C70EC",
x"8F18723E",
x"9056734B",
x"913F73F8",
x"91C6743B",
x"91ED7412",
x"91BB738B",
x"914272B9",
x"90A171BB",
x"8FF270B1",
x"8F566FB3",
x"8EE66ED7",
x"8EB26E2A",
x"8EC16DB0",
x"8F0E6D65",
x"8F8B6D44",
x"90256D3F",
x"90C16D51",
x"91496D6F",
x"91AB6D99",
x"91D96DCA",
x"91D26E06",
x"91986E4A",
x"91366E96",
x"90B86EE4",
x"902C6F2D",
x"8FA26F69",
x"8F1F6F8D",
x"8EAE6F93",
x"8E4B6F78",
x"8DF66F3A",
x"8DAA6EDF",
x"8D606E72",
x"8D126DFC",
x"8CB86D89",
x"8C4B6D21",
x"8BC46CCB",
x"8B1B6C83",
x"8A4F6C48",
x"895A6C13",
x"88426BD9",
x"870E6B97",
x"85CF6B49",
x"849B6AF2",
x"838E6A96",
x"82C86A42",
x"82656A03",
x"827C69E5",
x"831B69F2",
x"84426A30",
x"85DC6A9C",
x"87C96B31",
x"89DF6BE1",
x"8BEA6C9D",
x"8DB86D52",
x"8F216DF3",
x"90086E73",
x"90626EC8",
x"90326EEF",
x"8F8D6EE5",
x"8E906EAE",
x"8D566E4D",
x"8BFB6DBF",
x"8A8E6D09",
x"89116C27",
x"87796B17",
x"85B169D5",
x"83A26863",
x"813B66C5",
x"7E6F6503",
x"7B45632D",
x"77D86156",
x"74515F97",
x"70E55E06",
x"6DD15CB9",
x"6B4B5BC3",
x"69805B2E",
x"68875AFA",
x"68665B24",
x"69095B9E",
x"6A485C57",
x"6BF05D3B",
x"6DCC5E33",
x"6FA75F31",
x"71566025",
x"72C46107",
x"73E661D3",
x"74C86289",
x"757C632D",
x"762163C4",
x"76D66456",
x"77B764EA",
x"78D56584",
x"7A376627",
x"7BDC66D3",
x"7DB4678A",
x"7FAC6848",
x"81AD6909",
x"839A69C8",
x"855F6A80",
x"86E96B2A",
x"882B6BC4",
x"89226C48",
x"89D06CB7",
x"8A3C6D13",
x"8A766D5F",
x"8A8E6DA3",
x"8A9B6DE8",
x"8AB26E37",
x"8AE66E96",
x"8B496F0C",
x"8BE76F9A",
x"8CC8703B",
x"8DE770EC",
x"8F4171A1",
x"90C87252",
x"926D72F2",
x"941E737E",
x"95C973EF",
x"9760744A",
x"98DA7492",
x"9A3174D1",
x"9B617512",
x"9C71755C",
x"9D6475B9",
x"9E407629",
x"9F0F76AD",
x"9FD67741",
x"A09777DB",
x"A1577877",
x"A217790C",
x"A2D57995",
x"A3927A0F",
x"A4497A7E",
x"A4F77AE5",
x"A5977B49",
x"A6227BAD",
x"A6917C16",
x"A6DD7C81",
x"A7017CED",
x"A6FA7D51",
x"A6C87DA8",
x"A6707DE7",
x"A5FD7E09",
x"A5787E0B",
x"A4F47DED",
x"A47E7DB2",
x"A4247D60",
x"A3ED7D02",
x"A3DC7CA0",
x"A3ED7C44",
x"A4177BF7",
x"A44C7BBA",
x"A47B7B91",
x"A4977B78",
x"A4917B6A",
x"A4637B5E",
x"A4087B4B",
x"A3877B29",
x"A2E67AEE",
x"A2307A92",
x"A1737A13",
x"A0B6796F",
x"A00178A7",
x"9F5477C0",
x"9EAE76C1",
x"9E0475B4",
x"9D4C74A0",
x"9C7E7392",
x"9B91728F",
x"9A8171A1",
x"995070CE",
x"9803701A",
x"96A76F86",
x"954B6F14",
x"93FE6EC5",
x"92CF6E96",
x"91C66E82",
x"90E76E86",
x"90326E9A",
x"8F9B6EB5",
x"8F176ECE",
x"8E9A6ED8",
x"8E146ECB",
x"8D816EA0",
x"8CDD6E51",
x"8C2F6DE2",
x"8B836D58",
x"8AE66CBD",
x"8A676C1E",
x"8A106B8C",
x"89E06B11",
x"89D06AB5",
x"89C86A7C",
x"89A76A5E",
x"89486A52",
x"88816A45",
x"872F6A24",
x"853C69DC",
x"82A1695C",
x"7F67689A",
x"7BAF6793",
x"77AB664E",
x"739464D5",
x"6FAD633F",
x"6C3161A1",
x"69556014",
x"673D5EAF",
x"65F95D86",
x"65845CA4",
x"65CB5C15",
x"66AA5BD7",
x"67F95BE9",
x"698A5C3F",
x"6B3A5CCD",
x"6CE65D86",
x"6E805E56",
x"6FFD5F33",
x"71636011",
x"72BD60E6",
x"741A61AF",
x"758C626C",
x"7721631E",
x"78E363CE",
x"7AD56481",
x"7CF3653F",
x"7F30660B",
x"817D66E9",
x"83C467D3",
x"85F068C7",
x"87ED69B8",
x"89A86A9D",
x"8B156B69",
x"8C2E6C12",
x"8CF16C8C",
x"8D656CD7",
x"8D926CF0",
x"8D8A6CDF",
x"8D5B6CAA",
x"8D186C5E",
x"8CD06C09",
x"8C936BB8",
x"8C656B79",
x"8C4C6B52",
x"8C486B4B",
x"8C566B62",
x"8C716B96",
x"8C916BDF",
x"8CAE6C34",
x"8CC26C8A",
x"8CC96CD7",
x"8CC16D10",
x"8CA56D31",
x"8C7A6D35",
x"8C3F6D1E",
x"8BF76CEF",
x"8BA56CAD",
x"8B4F6C5E",
x"8AF96C0A",
x"8AA56BB7",
x"8A5A6B69",
x"8A1A6B26",
x"89E76AEF",
x"89C36AC7",
x"89AD6AB0",
x"899F6AAD",
x"89976AC4",
x"898E6AF7",
x"897E6B4B",
x"89636BC4",
x"89396C62",
x"89006D20",
x"88BB6DF6",
x"88726EDB",
x"882E6FBE",
x"87F7708F",
x"87DB713E",
x"87E071BD",
x"880B7202",
x"885D7208",
x"88D371CF",
x"8963715F",
x"8A0170C3",
x"8AA17005",
x"8B356F35",
x"8BB16E65",
x"8C0D6D9E",
x"8C486CF0",
x"8C606C62",
x"8C5A6BFA",
x"8C406BBB",
x"8C186BA6",
x"8BE96BB7",
x"8BB56BE8",
x"8B806C31",
x"8B446C89",
x"8AFB6CE1",
x"8A9E6D2B",
x"8A246D5E",
x"89866D6E",
x"88BE6D52",
x"87D06D0C",
x"86C26C9C",
x"859D6C0C",
x"84706B68",
x"834C6ABD",
x"82416A1C",
x"815B6990",
x"80A46926",
x"801E68E2",
x"7FC968C7",
x"7F9D68CF",
x"7F9068F5",
x"7F946930",
x"7F9D6973",
x"7F9E69BA",
x"7F9069FA",
x"7F6A6A30",
x"7F286A56",
x"7ECB6A6B",
x"7E4F6A6B",
x"7DB26A51",
x"7CF36A16",
x"7C0D69B1",
x"7AF9691A",
x"79B26845",
x"78386731",
x"768965DE",
x"74A86450",
x"72A3629A",
x"708960CF",
x"6E6C5F0B",
x"6C665D6C",
x"6A8D5C0D",
x"68F75B05",
x"67BA5A64",
x"66DF5A2E",
x"66725A60",
x"66785AED",
x"66F25BC2",
x"67E25CCC",
x"69485DF6",
x"6B265F35",
x"6D7A6081",
x"704C61DD",
x"7397634F",
x"775964E2",
x"7B8766A3",
x"800D6897",
x"84D36AC2",
x"89B46D19",
x"8E8A6F8F",
x"932A720A",
x"976D7474",
x"9B2E76AD",
x"9E5678A2",
x"A0D77A3E",
x"A2B27B81",
x"A3F47C68",
x"A4B27D01",
x"A50F7D5B",
x"A52C7D91",
x"A52C7DB2",
x"A52B7DD1",
x"A5407DFA",
x"A5767E32",
x"A5CA7E77",
x"A6357EBF",
x"A6A27EFF",
x"A6FA7F2F",
x"A7257F40",
x"A70D7F2C",
x"A6A27EF2",
x"A5E07E95",
x"A4C97E1C",
x"A36E7D94",
x"A1E47D08",
x"A0467C89",
x"9EB37C1F",
x"9D457BCE",
x"9C117B99",
x"9B247B79",
x"9A817B65",
x"9A257B50",
x"9A057B2C",
x"9A107AEF",
x"9A347A93",
x"9A647A15",
x"9A947978",
x"9ABC78C7",
x"9AD9780F",
x"9AEA7760",
x"9AF376C4",
x"9AF3764B",
x"9AED75F8",
x"9AE075CB",
x"9ACC75C0",
x"9AAF75CB",
x"9A8875E4",
x"9A5A75F9",
x"9A297606",
x"99FB7602",
x"99D775EE",
x"99C375CD",
x"99C875A6",
x"99E37586",
x"9A147578",
x"9A577586",
x"9AA475B7",
x"9AF3760D",
x"9B3E7688",
x"9B847723",
x"9BC877D8",
x"9C10789C",
x"9C677965",
x"9CDC7A2F",
x"9D787AEF",
x"9E427BA5",
x"9F387C4A",
x"A0507CDB",
x"A1777D59",
x"A2957DB9",
x"A38C7DFA",
x"A43D7E12",
x"A48E7DFC",
x"A46E7DB0",
x"A3D67D2D",
x"A2CA7C72",
x"A15A7B88",
x"9FA47A77",
x"9DC3794E",
x"9BE07823",
x"9A177705",
x"98847602",
x"97397526",
x"963B7471",
x"958473DF",
x"95037365",
x"949E72F1",
x"9436726E",
x"93AC71CD",
x"92E37100",
x"91C57000",
x"90456ED2",
x"8E656D7F",
x"8C2F6C17",
x"89B96AB1",
x"87226961",
x"848D6838",
x"82156744",
x"7FD96687",
x"7DE665FF",
x"7C41659E",
x"7ADE6553",
x"79A16509",
x"786B64A5",
x"77106415",
x"756A6348",
x"73596232",
x"70C960D2",
x"6DB85F2C",
x"6A375D4D",
x"66635B49",
x"62725936",
x"5E995732",
x"5B155554",
x"581953BA",
x"55D25277",
x"545C519C",
x"53BE5132",
x"53EF5137",
x"54D751A8",
x"56525275",
x"5834538B",
x"5A5454D3",
x"5C895635",
x"5EB1579C",
x"60B858F7",
x"62905A39",
x"64355B5C",
x"65AB5C5F",
x"66FA5D46",
x"682D5E17",
x"69515EDA",
x"6A6D5F98",
x"6B8C6050",
x"6CB06107",
x"6DD961B8",
x"6F096259",
x"703862E3",
x"71636349",
x"727F6386",
x"73846390",
x"746A6366",
x"7528630B",
x"75B8628D",
x"761961F6",
x"764A6159",
x"765260CB",
x"763A605D",
x"760F6021",
x"75DE601E",
x"75B2605A",
x"759B60D3",
x"759E6181",
x"75BC6256",
x"75F66341",
x"76426431",
x"76976513",
x"76EB65D8",
x"77326673",
x"776966DC",
x"7787670E",
x"77916706",
x"778A66C8",
x"777D6655",
x"777065B7",
x"777264F3",
x"77866418",
x"77B46331",
x"77FA624C",
x"78596179",
x"78C960C8",
x"79456046",
x"79C56001",
x"7A446001",
x"7ABE6049",
x"7B3560D6",
x"7BAB619E",
x"7C236295",
x"7CA163A7",
x"7D2864BE",
x"7DB565C5",
x"7E4566A8",
x"7ECE675B",
x"7F4467D1",
x"7F976809",
x"7FBC6806",
x"7FA867D1",
x"7F556776",
x"7EC56704",
x"7DFF6689",
x"7D106610",
x"7C0D65A1",
x"7B096544",
x"7A1864F9",
x"794C64C1",
x"78B1649A",
x"78486481",
x"78136479",
x"7806647D",
x"7818648E",
x"783A64AA",
x"785D64CF",
x"787764F9",
x"78806521",
x"7872653C",
x"784E6542",
x"7814652B",
x"77C964EF",
x"7772648A",
x"77146401",
x"76B4635D",
x"765862AB",
x"76046200",
x"75C1616C",
x"75916104",
x"757A60D5",
x"758160E7",
x"75A5613B",
x"75E361C8",
x"7637627D",
x"76946346",
x"76F0640D",
x"773F64BB",
x"77776541",
x"77966590",
x"779865A7",
x"77876589",
x"776C6542",
x"775664DF",
x"77526470",
x"77656404",
x"779063A3",
x"77C6634E",
x"77F36300",
x"77F662AF",
x"77A8624B",
x"76E961C1",
x"75946103",
x"739A6007",
x"70F75ECC",
x"6DBE5D59",
x"6A165BC0",
x"66335A1B",
x"625B5887",
x"5ED45724",
x"5BE5560F",
x"59C55563",
x"589F552C",
x"58825570",
x"5969562B",
x"5B3A574D",
x"5DC858C2",
x"60DC5A73",
x"643E5C42",
x"67B15E1A",
x"6B075FE0",
x"6E1D6183",
x"70DB62F6",
x"7337642D",
x"75346525",
x"76DB65DC",
x"78376655",
x"79536696",
x"7A3E66AA",
x"7AFD669A",
x"7B966673",
x"7C0D6642",
x"7C686614",
x"7CAA65F0",
x"7CDE65DE",
x"7D0B65DF",
x"7D4165F2",
x"7D876610",
x"7DE96632",
x"7E696652",
x"7F046668",
x"7FB5666D",
x"806D6665",
x"811E664E",
x"81B7662E",
x"822B660E",
x"827265F5",
x"828665E9",
x"826965F0",
x"8227660A",
x"81C56635",
x"8155666F",
x"80E266B0",
x"807666F3",
x"801A6735",
x"7FD66772",
x"7FAF67AB",
x"7FA867E3",
x"7FC56823",
x"8009686C",
x"807668C5",
x"810E6931",
x"81CE69B0",
x"82AF6A3D",
x"83A86AD1",
x"84A76B65",
x"85976BED",
x"86636C65",
x"86FA6CC1",
x"87496CFF",
x"874B6D21",
x"87016D2A",
x"867A6D20",
x"85CC6D0C",
x"85136CF6",
x"846C6CE9",
x"83F66CE9",
x"83C26CF9",
x"83DD6D1C",
x"84446D4D",
x"84E66D89",
x"85AB6DC8",
x"86746E03",
x"87216E34",
x"87926E54",
x"87B56E5E",
x"87806E4F",
x"86F76E29",
x"86286DE9",
x"852F6D96",
x"84286D34",
x"83326CC7",
x"82656C57",
x"81D26BE6",
x"817D6B7C",
x"81626B1C",
x"816D6AC8",
x"818B6A82",
x"81A26A49",
x"81976A20",
x"81596A00",
x"80DC69E9",
x"802069D6",
x"7F2C69C4",
x"7E1169AB",
x"7CE26989",
x"7BB76959",
x"7AA3691B",
x"79BA68CE",
x"79046875",
x"788D6816",
x"784F67B7",
x"78486760",
x"786C671A",
x"78B266EB",
x"791066D8",
x"797966E0",
x"79E96706",
x"7A5B6741",
x"7ACE678A",
x"7B4167D9",
x"7BB76824",
x"7C2E6862",
x"7CA5688C",
x"7D176899",
x"7D776886",
x"7DB76851",
x"7DC567F6",
x"7D936777",
x"7D1366D9",
x"7C3F661E",
x"7B1D6553",
x"79BC6486",
x"783B63C5",
x"76C26325",
x"758362BE",
x"74AF62A1",
x"747962DD",
x"7507637F",
x"76726486",
x"78C165E9",
x"7BE96799",
x"7FCF697D",
x"84486B7F",
x"891F6D85",
x"8E1E6F76",
x"9311714A",
x"97CC72F8",
x"9C2B7485",
x"A01C75FC",
x"A398776F",
x"A6A578EE",
x"A9507A89",
x"ABB37C4D",
x"ADE37E3A",
x"AFFD804F",
x"B2168282",
x"B43D84C3",
x"B67B86FD",
x"B8CF891D",
x"BB2D8B0E",
x"BD898CC2",
x"BFCC8E2C",
x"C1DE8F4B",
x"C3AA901B",
x"C52290A5",
x"C63C90F3",
x"C6FB9113",
x"C76A9116",
x"C79C910C",
x"C7AB9103",
x"C7B09107",
x"C7CC911E",
x"C80E9148",
x"C889917F",
x"C94391B8",
x"CA3A91E9",
x"CB689202",
x"CCC091FC",
x"CE3791D3",
x"CFC3918D",
x"D15B9134",
x"D2F990DD",
x"D49F90A1",
x"D64B9097",
x"D80290D3",
x"D9C19166",
x"DB89924E",
x"DD549384",
x"DF1994F2",
x"E0CE967C",
x"E26797FC",
x"E3D09952",
x"E4FB9A61",
x"E5D89B15",
x"E65E9B62",
x"E6809B51",
x"E63E9AF1",
x"E5999A5A",
x"E49D99A7",
x"E35B98F9",
x"E1EB9868",
x"E06C9803",
x"DEFC97D2",
x"DDBC97D5",
x"DCC19800",
x"DC1F9844",
x"DBDA988F",
x"DBEC98CE",
x"DC4698F9",
x"DCCE9909",
x"DD689900",
x"DDF998E8",
x"DE6998CC",
x"DEAA98BB",
x"DEB898C4",
x"DE9998EF",
x"DE579940",
x"DE0299B3",
x"DDA79A3D",
x"DD529ACE",
x"DD089B55",
x"DCC09BC1",
x"DC749C06",
x"DC169C1C",
x"DB989C00",
x"DAF49BBD",
x"DA249B5B",
x"D9349AE6",
x"D8339A6C",
x"D73199F6",
x"D6489989",
x"D58B9920",
x"D50898B8",
x"D4C69848",
x"D4C397C8",
x"D4F69733",
x"D554968A",
x"D5CB95D5",
x"D6509524",
x"D6DA948A",
x"D7649420",
x"D7EF93F6",
x"D87C941A",
x"D90F9490",
x"D9A49552",
x"DA3A964A",
x"DAC79760",
x"DB409876",
x"DB96996E",
x"DBC39A2D",
x"DBBD9AA3",
x"DB7F9ACB",
x"DB099AA4",
x"DA589A3A",
x"D9679991",
x"D82698B5",
x"D68297A4",
x"D4589656",
x"D18194BB",
x"CDD392B9",
x"C92A9039",
x"C3758D27",
x"BCB8897A",
x"B512853F",
x"ACC78092",
x"A4327BA8",
x"9BC276C1",
x"93F17229",
x"8D346E2D",
x"87EA6B10",
x"84566900",
x"82976819",
x"82A36858",
x"844969A0",
x"87436BC2",
x"8B386E80",
x"8FCB719C",
x"94A874D5",
x"998A77FB",
x"9E457AEE",
x"A2BF7D9C",
x"A6F58005",
x"AAF18239",
x"AEBF8443",
x"B2708636",
x"B60E881F",
x"B99889FE",
x"BD088BD0",
x"C04E8D8B",
x"C35A8F1B",
x"C61B9074",
x"C885918D",
x"CA93925D",
x"CC4992F0",
x"CDAF934F",
x"CED4938D",
x"CFC893BF",
x"D09B93F6",
x"D155943F",
x"D1FE949E",
x"D292950A",
x"D30C9579",
x"D36295D8",
x"D38E9614",
x"D382961E",
x"D33A95EE",
x"D2B29582",
x"D1EB94E0",
x"D0E89417",
x"CFB3933B",
x"CE54925F",
x"CCDB9197",
x"CB5590F3",
x"C9D8907D",
x"C878903C",
x"C74E9035",
x"C6749067",
x"C60290D2",
x"C6109172",
x"C6AD9245",
x"C7E09349",
x"C99D9476",
x"CBD495C4",
x"CE609724",
x"D1109885",
x"D3B699CF",
x"D6199AF3",
x"D80C9BDC",
x"D96F9C80",
x"DA319CD8",
x"DA559CE8",
x"D9EE9CBA",
x"D91F9C5B",
x"D8139BDF",
x"D6F99B54",
x"D5FB9ACA",
x"D5399A45",
x"D4C799CC",
x"D4A7995F",
x"D4D498FB",
x"D53B989F",
x"D5C6984E",
x"D65E980D",
x"D6EF97E5",
x"D77197DF",
x"D7DB9803",
x"D8339854",
x"D88198CC",
x"D8CE995E",
x"D92499F8",
x"D98F9A80",
x"DA0C9AE4",
x"DA9D9B0D",
x"DB3E9AF8",
x"DBEA9AA7",
x"DC969A2B",
x"DD40999F",
x"DDE49923",
x"DE8598DA",
x"DF2498DF",
x"DFC79944",
x"E0719A0A",
x"E1239B29",
x"E1DD9C83",
x"E2939DF5",
x"E3399F52",
x"E3BBA075",
x"E403A139",
x"E3F6A185",
x"E380A14B",
x"E28CA08F",
x"E10C9F5B",
x"DEFC9DC4",
x"DC619BE4",
x"D94A99D5",
x"D5CA97B4",
x"D1FF9594",
x"CE099389",
x"CA07919A",
x"C6168FD1",
x"C2518E2B",
x"BECD8CA8",
x"BB958B42",
x"B8AF89F1",
x"B61888AC",
x"B3C28767",
x"B1968615",
x"AF7884A9",
x"AD408311",
x"AAC3813B",
x"A7CF7F18",
x"A4387C9B",
x"9FDA79B9",
x"9AA17672",
x"948672CD",
x"8DA06EDE",
x"861B6AC2",
x"7E4266A1",
x"766962A7",
x"6EF65F07",
x"684F5BF0",
x"62CC5988",
x"5EB857ED",
x"5C3D5729",
x"5B62573A",
x"5C14580A",
x"5E1E5971",
x"61355B45",
x"65025D4F",
x"692A5F5F",
x"6D596149",
x"714C62EF",
x"74D4643C",
x"77D26532",
x"7A4265D8",
x"7C2F6642",
x"7DB4668B",
x"7EED66D1",
x"8000672A",
x"810C67AA",
x"822A685E",
x"836F6947",
x"84E56A5F",
x"868B6B9C",
x"885F6CEC",
x"8A506E3E",
x"8C4F6F7F",
x"8E4370A0",
x"901A7196",
x"91C2725B",
x"932E72EF",
x"94577358",
x"953F73A0",
x"95EA73D5",
x"96667405",
x"96BD743B",
x"97017483",
x"973974E1",
x"976E7555",
x"97A175D8",
x"97D27660",
x"97FB76DB",
x"981D773C",
x"98367775",
x"984A777E",
x"98637755",
x"988D7702",
x"98D6768F",
x"994C7612",
x"99F7759C",
x"9ADC7544",
x"9BF1751C",
x"9D2E752D",
x"9E7A757B",
x"9FC27602",
x"A0F076B4",
x"A1F07781",
x"A2B87854",
x"A349791C",
x"A3AC79C9",
x"A3F67A56",
x"A4407AC1",
x"A4AE7B1C",
x"A5607B77",
x"A6787BEE",
x"A80F7CA0",
x"AA3B7DAA",
x"ACFE7F25",
x"B056811F",
x"B430839E",
x"B86E8691",
x"BCE489E2",
x"C1608D67",
x"C5AA90F2",
x"C98F944E",
x"CCE1974A",
x"CF7E99BA",
x"D1539B82",
x"D25E9C95",
x"D2AF9CF6",
x"D25F9CBB",
x"D1969C02",
x"D07E9AF2",
x"CF3A99B3",
x"CDE89868",
x"CC9D972B",
x"CB5F960D",
x"CA29950D",
x"C8EE9424",
x"C79D9342",
x"C6289256",
x"C485914E",
x"C2B3901E",
x"C0BC8EC5",
x"BEB08D48",
x"BCA88BB5",
x"BABF8A24",
x"B90F88AB",
x"B7B38766",
x"B6BD866D",
x"B63585CF",
x"B61F8597",
x"B67385C6",
x"B7238656",
x"B81C8735",
x"B944884C",
x"BA7E8980",
x"BBA98AB2",
x"BCA88BC3",
x"BD608C9B",
x"BDB78D24",
x"BD9F8D4E",
x"BD118D14",
x"BC0C8C79",
x"BA978B84",
x"B8BC8A42",
x"B68B88C0",
x"B40B870D",
x"B142852F",
x"AE2E832C",
x"AAC98102",
x"A70A7EB2",
x"A2E77C32",
x"9E637983",
x"998876AC",
x"947373BA",
x"8F5070C4",
x"8A5C6DE8",
x"85D96B4B",
x"820D6911",
x"7F346758",
x"7D796637",
x"7CF065B7",
x"7D8E65D3",
x"7F30667C",
x"819B6791",
x"848968F3",
x"87AC6A7D",
x"8AC26C14",
x"8D976DA3",
x"900E6F21",
x"92257093",
x"93EA7206",
x"9583738C",
x"97177539",
x"98D2771C",
x"9AD6793D",
x"9D387B9B",
x"9FFB7E23",
x"A31580C3",
x"A66A835D",
x"A9DA85D3",
x"AD40880A",
x"B07D89EA",
x"B3748B69",
x"B6128C80",
x"B84D8D36",
x"BA228D98",
x"BB938DB6",
x"BCAC8DA4",
x"BD748D74",
x"BDFB8D3B",
x"BE4F8D08",
x"BE848CE9",
x"BEAF8CE7",
x"BEEA8D0D",
x"BF4A8D5B",
x"BFEA8DD2",
x"C0D68E6D",
x"C2188F21",
x"C3B08FE3",
x"C58E90A1",
x"C796914B",
x"C9AA91D2",
x"CBA3922E",
x"CD5D925B",
x"CEBD925C",
x"CFB69244",
x"D04A9223",
x"D08C9213",
x"D09F922D",
x"D0AC9284",
x"D0E49327",
x"D16E9416",
x"D2659548",
x"D3D896AA",
x"D5BD9820",
x"D7F7998D",
x"DA5E9AD4",
x"DCBE9BDC",
x"DEE79C96",
x"E0AD9CFC",
x"E1F29D0C",
x"E2AF9CD4",
x"E2E89C5C",
x"E2B99BB6",
x"E2449AEC",
x"E1B39A06",
x"E12A9909",
x"E0C197F5",
x"E08596C5",
x"E06F957C",
x"E06E9417",
x"E05F929E",
x"E020911A",
x"DF8F8F9B",
x"DE928E32",
x"DD198CF3",
x"DB258BEA",
x"D8C18B24",
x"D6058AA4",
x"D30E8A66",
x"CFF48A5C",
x"CCD48A74",
x"C9BD8A9B",
x"C6B98AB8",
x"C3CC8AB5",
x"C0F28A81",
x"BE2D8A10",
x"BB78895C",
x"B8DB8866",
x"B65B8733",
x"B40785CC",
x"B1EB843F",
x"B016829B",
x"AE9280F0",
x"AD607F4D",
x"AC7B7DC4",
x"ABD67C64",
x"AB5D7B3C",
x"AAFD7A57",
x"AA9E79C0",
x"AA2F7979",
x"A9A47982",
x"A8F179D1",
x"A8177A56",
x"A7147AF9",
x"A5EB7BA0",
x"A4A17C2D",
x"A3387C84",
x"A1B57C8C",
x"A0197C37",
x"9E6A7B7F",
x"9CAC7A68",
x"9AE97902",
x"99287767",
x"977375AF",
x"95CD73F5",
x"943B7254",
x"92B670D7",
x"91316F82",
x"8F9A6E4F",
x"8DD66D31",
x"8BD26C13",
x"89766AE1",
x"86B8698A",
x"839F680A",
x"80396660",
x"7CAB649E",
x"792062D9",
x"75CC6131",
x"72E65FC5",
x"709B5EB1",
x"6F105E0A",
x"6E595DD9",
x"6E785E1C",
x"6F5B5EC8",
x"70E85FC6",
x"72F760FA",
x"7560624C",
x"77FA63A4",
x"7AA164F0",
x"7D3C6627",
x"7FBB6744",
x"8210684B",
x"843C6944",
x"86416A32",
x"881D6B1D",
x"89D36C09",
x"8B666CF5",
x"8CD06DDF",
x"8E116EC3",
x"8F256F9C",
x"900D7065",
x"90C9711D",
x"916271C1",
x"91DC7254",
x"924572D4",
x"92A77343",
x"931073A3",
x"938B73F6",
x"9421743D",
x"94DC7479",
x"95BF74B1",
x"96D374EA",
x"981B752C",
x"99977582",
x"9B4B75F9",
x"9D31769C",
x"9F497774",
x"A1887888",
x"A3E779DB",
x"A6547B67",
x"A8C07D20",
x"AB187EFB",
x"AD4880DE",
x"AF4082B6",
x"B0F08467",
x"B24D85DA",
x"B35086FA",
x"B3F787B6",
x"B4428808",
x"B43887EE",
x"B3E48773",
x"B35386A7",
x"B294859F",
x"B1B7847A",
x"B0D38354",
x"AFF58249",
x"AF328172",
x"AE9B80E1",
x"AE3F809F",
x"AE2B80AF",
x"AE69810A",
x"AEFF81A3",
x"AFF0826E",
x"B1388359",
x"B2D18453",
x"B4B08552",
x"B6C2864A",
x"B8F28738",
x"BB2B8817",
x"BD4C88E4",
x"BF39899D",
x"C0D88A3E",
x"C20E8AC0",
x"C2C68B1E",
x"C2F58B4F",
x"C2988B4B",
x"C1B78B11",
x"C0678AA2",
x"BEC18A07",
x"BCEA894A",
x"BB09887B",
x"B94487AF",
x"B7BD86F6",
x"B68F865E",
x"B5C685F0",
x"B56485AE",
x"B5608592",
x"B5A38592",
x"B611859E",
x"B68485A5",
x"B6DA8597",
x"B6F48566",
x"B6B8850D",
x"B619848B",
x"B51883E6",
x"B3BC8328",
x"B21E8260",
x"B05D819F",
x"AE9C80F7",
x"AD078075",
x"ABBB8026",
x"AAD48012",
x"AA66803D",
x"AA7180A5",
x"AAED8142",
x"ABC2820A",
x"ACCF82EB",
x"ADF083D6",
x"AF0184B2",
x"AFE4856E",
x"B08785F8",
x"B0E18640",
x"B0FA863D",
x"B0DD85F0",
x"B0A18559",
x"B0538481",
x"AFFD8374",
x"AF99823C",
x"AF1180E1",
x"AE3C7F68",
x"ACE77DCF",
x"AAD77C09",
x"A7DC7A0F",
x"A3CD77D1",
x"9EA57547",
x"98747272",
x"91736F59",
x"89F76C14",
x"826A68C5",
x"7B456597",
x"74FC62B9",
x"6FF56059",
x"6C785E9B",
x"6AAA5D97",
x"6A865D53",
x"6BDF5DC1",
x"6E6F5EC1",
x"71D2602B",
x"75A161CC",
x"79776373",
x"7D0064F6",
x"7FFF6638",
x"8250672D",
x"83F067D3",
x"84F06841",
x"8576688D",
x"85AC68D5",
x"85C56937",
x"85E769C5",
x"86346A87",
x"86B96B7C",
x"877C6C92",
x"88706DB3",
x"89876EC4",
x"8AA76FAB",
x"8BB97057",
x"8CAC70B9",
x"8D7170D2",
x"8E0470AB",
x"8E667052",
x"8E9B6FD9",
x"8EAB6F54",
x"8E9F6ECE",
x"8E7E6E52",
x"8E486DDF",
x"8DFC6D73",
x"8D926D08",
x"8D066C92",
x"8C4F6C0F",
x"8B696B7D",
x"8A566AE3",
x"891F6A4C",
x"87D669C7",
x"86906962",
x"8566692D",
x"84746931",
x"83D06970",
x"838D69E8",
x"83AF6A8C",
x"84356B4E",
x"85146C21",
x"86356CF5",
x"87836DBF",
x"88E46E7F",
x"8A426F31",
x"8B8D6FDE",
x"8CBC708A",
x"8DCD7140",
x"8EC67200",
x"8FAB72CE",
x"908673A3",
x"91597475",
x"92247537",
x"92E075DA",
x"9381764E",
x"93F4768B",
x"942B7688",
x"94147647",
x"93A575CA",
x"92DF751C",
x"91C87448",
x"9071735E",
x"8EF9726B",
x"8D7E717E",
x"8C2570A3",
x"8B0E6FE5",
x"8A596F4D",
x"8A176EDF",
x"8A536EA3",
x"8B0B6E96",
x"8C2F6EB7",
x"8DA76F02",
x"8F526F6C",
x"910A6FE8",
x"92AB7069",
x"941070E1",
x"951C713D",
x"95BE7172",
x"95E97178",
x"959F714B",
x"94EC70EE",
x"93E57069",
x"92A16FCD",
x"91406F26",
x"8FDC6E89",
x"8E916E06",
x"8D736DA7",
x"8C8E6D78",
x"8BEC6D76",
x"8B896DA0",
x"8B5F6DEB",
x"8B656E48",
x"8B8A6EAA",
x"8BC06F05",
x"8BFB6F4D",
x"8C326F7A",
x"8C5C6F8D",
x"8C7B6F88",
x"8C946F70",
x"8CAB6F52",
x"8CCB6F35",
x"8CFB6F23",
x"8D426F21",
x"8D986F30",
x"8DF76F4A",
x"8E486F62",
x"8E706F68",
x"8E4D6F45",
x"8DBE6EE4",
x"8C9D6E2D",
x"8AD36D13",
x"88566B8F",
x"852B69A4",
x"816A675F",
x"7D3F64DE",
x"78E36241",
x"74965FB3",
x"709B5D60",
x"6D315B6E",
x"6A8959FD",
x"68C1591F",
x"67E658DD",
x"67EC592C",
x"68B759F7",
x"6A1D5B21",
x"6BEF5C86",
x"6DFA5E03",
x"70115F76",
x"721160C9",
x"73E561EF",
x"758362E0",
x"76ED63A7",
x"7832644C",
x"796264E5",
x"7A91657D",
x"7BD26628",
x"7D3166EF",
x"7EB567D3",
x"805F68D6",
x"822569ED",
x"83FC6B10",
x"85D36C2E",
x"879A6D3F",
x"893F6E38",
x"8AB66F13",
x"8BF96FCD",
x"8D07706B",
x"8DE570F0",
x"8E9E7169",
x"8F4171DB",
x"8FDD7250",
x"908472CB",
x"913E734E",
x"921573D5",
x"9307745C",
x"941074DA",
x"95217543",
x"962E7590",
x"972475BC",
x"97F475C1",
x"989475A3",
x"98FE756B",
x"9934751F",
x"993C74D0",
x"9925748B",
x"9900745B",
x"98DA744A",
x"98C6745C",
x"98CA7492",
x"98EE74E4",
x"9932754A",
x"999575B9",
x"9A117625",
x"9AA17686",
x"9B4076D5",
x"9BEA7713",
x"9C9C7741",
x"9D557764",
x"9E0E7782",
x"9EC677A3",
x"9F7477CE",
x"A00E7803",
x"A0887843",
x"A0DA7889",
x"A0FB78D0",
x"A0EB7910",
x"A0AC7943",
x"A0497962",
x"9FD2796B",
x"9F57795D",
x"9EED7937",
x"9EA478FF",
x"9E8478BC",
x"9E94786F",
x"9ECD7822",
x"9F2777D7",
x"9F8E778F",
x"9FF4774E",
x"A0467712",
x"A07976D8",
x"A080769F",
x"A05A7662",
x"A0087623",
x"9F8F75DB",
x"9EF1758D",
x"9E337539",
x"9D5774DC",
x"9C5D747C",
x"9B437419",
x"9A0573B6",
x"98A47355",
x"972172F8",
x"958172A0",
x"93D2724B",
x"921D71F8",
x"907471A3",
x"8EE97147",
x"8D8770DF",
x"8C597066",
x"8B636FD9",
x"8AA26F38",
x"8A136E86",
x"89A86DCA",
x"89566D0A",
x"89116C54",
x"88CE6BB4",
x"88836B34",
x"882E6ADF",
x"87CF6ABA",
x"87666AC4",
x"86F96AF6",
x"86886B47",
x"86186BA6",
x"85A56BFF",
x"852C6C3E",
x"84A86C51",
x"840E6C27",
x"83586BB4",
x"827A6AF6",
x"817269EF",
x"803868AA",
x"7ED36735",
x"7D4865A7",
x"7BA36415",
x"79F3629A",
x"784E6148",
x"76C46031",
x"756A5F60",
x"74535EDD",
x"738C5EA8",
x"731D5EB9",
x"73095F06",
x"734F5F83",
x"73E8601E",
x"74C860CC",
x"75E26183",
x"7727623B",
x"788C62EF",
x"7A0363A1",
x"7B8A6456",
x"7D1E6514",
x"7EBF65E2",
x"807366C4",
x"823E67BC",
x"842068CE",
x"861869F6",
x"88226B2D",
x"8A346C6C",
x"8C3F6DAA",
x"8E346EDE",
x"90037002",
x"91A1710F",
x"93077200",
x"943572D7",
x"95327390",
x"96067431",
x"96BF74BA",
x"976D752F",
x"981E7592",
x"98D875E8",
x"999F7634",
x"9A76767E",
x"9B5376C7",
x"9C327716",
x"9D0A7771",
x"9DD577DB",
x"9E8E7856",
x"9F3578E1",
x"9FCD7977",
x"A05A7A12",
x"A0E37AA9",
x"A16D7B32",
x"A2017BA6",
x"A2A17BFE",
x"A3527C39",
x"A4177C59",
x"A4F47C65",
x"A5EB7C68",
x"A6FD7C6F",
x"A8287C85",
x"A9677CB3",
x"AAB37CFC",
x"AC007D61",
x"AD397DD7",
x"AE4D7E54",
x"AF267EC6",
x"AFB27F1F",
x"AFE07F50",
x"AFAB7F50",
x"AF157F1C",
x"AE2E7EBA",
x"AD0B7E2F",
x"ABC97D8E",
x"AA887CE7",
x"A96B7C50",
x"A88E7BD7",
x"A8057B89",
x"A7DD7B6F",
x"A8177B86",
x"A8AB7BCD",
x"A98B7C39",
x"AAA67CBD",
x"ABE87D4E",
x"AD3D7DE0",
x"AE997E65",
x"AFEE7EDA",
x"B1357F37",
x"B26A7F81",
x"B3897FB6",
x"B4927FDB",
x"B5827FF7",
x"B656800F",
x"B707802B",
x"B791804A",
x"B7EB8070",
x"B811809B",
x"B7F780C6",
x"B79680EA",
x"B6E880FA",
x"B5E780ED",
x"B48C80B7",
x"B2D7804D",
x"B0C77FAB",
x"AE637ECD",
x"ABB27DB6",
x"A8C57C72",
x"A5B27B0E",
x"A29579A0",
x"9F8E783E",
x"9CBD76FE",
x"9A4075F1",
x"982F7527",
x"969774A6",
x"95797468",
x"94C87465",
x"946D7488",
x"944874B9",
x"943474DE",
x"940D74E1",
x"93B574AC",
x"931A7437",
x"9235737E",
x"910E7288",
x"8FB57161",
x"8E45701F",
x"8CD36ED5",
x"8B796D96",
x"8A3B6C6C",
x"891B6B5F",
x"88066A69",
x"86DF6982",
x"85866896",
x"83D86796",
x"81B86670",
x"7F1B651A",
x"7C046393",
x"788E61E0",
x"74E56015",
x"713F5E4D",
x"6DDE5CA7",
x"6B005B40",
x"68DB5A36",
x"6790599E",
x"67315980",
x"67B359D9",
x"68FC5A9B",
x"6ADB5BB1",
x"6D1B5CF7",
x"6F835E50",
x"71D95F9B",
x"73F860BF",
x"75BE61A9",
x"77246253",
x"782B62C4",
x"78E66304",
x"796F632D",
x"79E36355",
x"7A636394",
x"7B0763FF",
x"7BE364A3",
x"7CFD6581",
x"7E56669A",
x"7FE567DB",
x"81976930",
x"83586A83",
x"85116BBB",
x"86AF6CC5",
x"88216D93",
x"895C6E21",
x"8A5F6E73",
x"8B2E6E96",
x"8BD56E9E",
x"8C636E9E",
x"8CED6EAE",
x"8D866EDE",
x"8E3C6F35",
x"8F1D6FB7",
x"902B705C",
x"91647116",
x"92C071D1",
x"942B7278",
x"959472F9",
x"96E27348",
x"9804735F",
x"98EA7343",
x"998D7302",
x"99ED72AD",
x"9A14725F",
x"9A147230",
x"9A087233",
x"9A0E7279",
x"9A3F730B",
x"9AB873E2",
x"9B8874F6",
x"9CB87634",
x"9E427788",
x"A01478D6",
x"A2147A09",
x"A41A7B0F",
x"A6017BDA",
x"A79E7C63",
x"A8D07CAC",
x"A97B7CB9",
x"A9927C96",
x"A9157C53",
x"A8127BF9",
x"A6A57B9B",
x"A4F07B41",
x"A31C7AF2",
x"A1577AB6",
x"9FC87A8B",
x"9E8E7A71",
x"9DC27A63",
x"9D717A5E",
x"9D9A7A61",
x"9E337A65",
x"9F2E7A6F",
x"A06E7A7F",
x"A1DA7A9B",
x"A3597AC9",
x"A4CF7B0C",
x"A6287B6F",
x"A7547BF2",
x"A8467C96",
x"A8F47D54",
x"A95B7E25",
x"A97A7EF8",
x"A94A7FBD",
x"A8D08064",
x"A80A80D7",
x"A6FD8108",
x"A5AC80ED",
x"A4218081",
x"A2667FC3",
x"A08B7EBD",
x"9EA27D7C",
x"9CBD7C11",
x"9AF17A8E",
x"994F7906",
x"97E97790",
x"96C6763A",
x"95EE750F",
x"955D7416",
x"950A7352",
x"94E472C1",
x"94D67258",
x"94C9720F",
x"94A471D7",
x"945271A1",
x"93C67162",
x"92F9710D",
x"91ED709D",
x"90B17010",
x"8F5A6F6C",
x"8E046EBB",
x"8CC96E0A",
x"8BBF6D6C",
x"8AF76CEB",
x"8A706C93",
x"8A1E6C66",
x"89E36C5F",
x"899A6C72",
x"89136C86",
x"88206C82",
x"86976C4A",
x"84636BC4",
x"817C6AE1",
x"7DF66996",
x"79F767E9",
x"75BB65EF",
x"718963C2",
x"6DAA618A",
x"6A655F6C",
x"67F35D92",
x"667C5C1B",
x"660C5B1C",
x"669E5AA1",
x"68145AA1",
x"6A425B10",
x"6CF25BD0",
x"6FE95CC8",
x"72F35DD9",
x"75E05EEC",
x"78915FEE",
x"7AF360DC",
x"7CFD61B8",
x"7EB7628D",
x"802D636A",
x"81706463",
x"829A6584",
x"83BC66D6",
x"84EA6858",
x"86316A03",
x"879B6BC5",
x"892D6D89",
x"8AE66F35",
x"8CC570B9",
x"8EC171FE",
x"90D572FC",
x"92F373B4",
x"95127430",
x"9727747E",
x"992474B4",
x"9AFD74EB",
x"9CA87536",
x"9E1C75A6",
x"9F537646",
x"A0497712",
x"A1037803",
x"A187790B",
x"A1E17A12",
x"A2257B04",
x"A2647BCE",
x"A2B37C64",
x"A3267CBF",
x"A3CA7CE1",
x"A4A87CD7",
x"A5BC7CB2",
x"A6FE7C89",
x"A8617C71",
x"A9D07C7E",
x"AB387CBC",
x"AC877D32",
x"ADAC7DDA",
x"AEA57EAD",
x"AF6E7F98",
x"B00C808B",
x"B0878170",
x"B0E68237",
x"B12D82D4",
x"B1608340",
x"B178837A",
x"B1728382",
x"B1498366",
x"B0F8832B",
x"B08582DE",
x"AFFB828C",
x"AF738242",
x"AF05820A",
x"AED781EE",
x"AF0581F7",
x"AFAB822B",
x"B0D3828F",
x"B27D8322",
x"B49283E1",
x"B6F184C5",
x"B96A85BF",
x"BBCC86C0",
x"BDE587B9",
x"BF8B8897",
x"C0A5894D",
x"C12689D3",
x"C1188A25",
x"C08F8A45",
x"BFAC8A3C",
x"BE948A17",
x"BD6A89E6",
x"BC4E89B5",
x"BB568991",
x"BA89897D",
x"B9EA897B",
x"B96D8983",
x"B9078988",
x"B8A58980",
x"B83D895A",
x"B7C3890B",
x"B736888E",
x"B69887E3",
x"B5F0870F",
x"B5448621",
x"B49E8527",
x"B3FE8433",
x"B3648356",
x"B2C58298",
x"B20E8200",
x"B12C8187",
x"B0088125",
x"AE9480C9",
x"ACC68061",
x"AA9E7FDB",
x"A82B7F2D",
x"A5877E4F",
x"A2D97D41",
x"A0457C11",
x"9DF37ACB",
x"9BFE7988",
x"9A797858",
x"995A774B",
x"9893766A",
x"97F775B1",
x"97597516",
x"96837485",
x"954673E5",
x"937E7320",
x"911F721F",
x"8E2B70D5",
x"8AC26F43",
x"87116D6E",
x"83556B70",
x"7FCB6966",
x"7CAF6776",
x"7A3465C5",
x"78796474",
x"778D639F",
x"77706358",
x"780E63A1",
x"79516474",
x"7B1865C1",
x"7D45676B",
x"7FC16958",
x"82766B69",
x"85566D82",
x"885A6F8D",
x"8B7D7179",
x"8EB87340",
x"920474DE",
x"95597658",
x"98AE77B7",
x"9BF47909",
x"9F247A57",
x"A2337BAA",
x"A51B7D09",
x"A7DC7E7A",
x"AA777FF7",
x"ACEE8180",
x"AF47830C",
x"B1888497",
x"B3B28615",
x"B5C38781",
x"B7B688D2",
x"B9848A00",
x"BB268B08",
x"BC948BE5",
x"BDC68C91",
x"BEBD8D0D",
x"BF7A8D59",
x"C0018D7A",
x"C05E8D74",
x"C09D8D56",
x"C0CC8D2B",
x"C0F58D01",
x"C1268CEA",
x"C1668CF3",
x"C1B68D27",
x"C2188D8A",
x"C2858E1E",
x"C2F88EDB",
x"C3688FB5",
x"C3D3909D",
x"C4329182",
x"C4899255",
x"C4E0930C",
x"C540939B",
x"C5BA9407",
x"C658944F",
x"C723947D",
x"C81C9499",
x"C93794A8",
x"CA6194B1",
x"CB7994B1",
x"CC5B94A5",
x"CCDE9486",
x"CCE49445",
x"CC5593DE",
x"CB309348",
x"C9859287",
x"C77B91A2",
x"C54690AB",
x"C3298FB9",
x"C1628EE7",
x"C02C8E53",
x"BFAB8E13",
x"BFEE8E35",
x"C0EA8EC1",
x"C2778FAF",
x"C45D90EA",
x"C6579258",
x"C81D93CF",
x"C9729528",
x"CA26963E",
x"CA2296EE",
x"C9649723",
x"C7FE96D1",
x"C61695FA",
x"C3D994AE",
x"C1779304",
x"BF1F911B",
x"BCF18F17",
x"BB088D18",
x"B96A8B3E",
x"B818899F",
x"B705884A",
x"B61F8748",
x"B554868F",
x"B48C8615",
x"B3B985C8",
x"B2CA858D",
x"B1B7854D",
x"B08084F1",
x"AF24846A",
x"ADA983AB",
x"AC1F82B3",
x"AA91818A",
x"A90C803F",
x"A7A27EE7",
x"A65D7D96",
x"A5467C68",
x"A4607B6F",
x"A3A97ABA",
x"A31F7A4D",
x"A2B67A2A",
x"A26B7A47",
x"A2367A96",
x"A2147B0B",
x"A2037B91",
x"A2037C18",
x"A2147C95",
x"A22C7CFA",
x"A23C7D39",
x"A2257D44",
x"A1BF7D0B",
x"A0D67C7B",
x"9F367B7F",
x"9CA87A03",
x"990777F7",
x"94427551",
x"8E65721A",
x"879E6E65",
x"803E6A58",
x"78AE6625",
x"716B620E",
x"6AF35E55",
x"65BF5B39",
x"622A58F4",
x"606F57A9",
x"60A0576B",
x"62A45833",
x"664459E7",
x"6B275C5D",
x"70EC5F5D",
x"772D62AF",
x"7D8E661D",
x"83C96977",
x"89A96C9D",
x"8F116F76",
x"93F471FB",
x"98547426",
x"9C3875FE",
x"9FA57788",
x"A29F78CD",
x"A52279D6",
x"A7297AA5",
x"A8AC7B43",
x"A9A67BB6",
x"AA1B7C04",
x"AA157C39",
x"A9A67C5E",
x"A8ED7C7F",
x"A80B7CA6",
x"A71F7CD7",
x"A6467D15",
x"A5947D5B",
x"A5127DA2",
x"A4C07DE0",
x"A4957E08",
x"A4817E11",
x"A4737DF2",
x"A4577DB0",
x"A4287D4D",
x"A3DF7CD6",
x"A3807C5A",
x"A3157BED",
x"A2AF7B9C",
x"A2597B75",
x"A2227B7E",
x"A2117BB9",
x"A2287C1C",
x"A2617C9F",
x"A2B37D30",
x"A3107DBF",
x"A3677E3C",
x"A3AB7E9C",
x"A3D37ED7",
x"A3DA7EEE",
x"A3BF7EE3",
x"A3877EBD",
x"A3397E87",
x"A2DF7E49",
x"A2807E0E",
x"A2227DD9",
x"A1C97DAA",
x"A1707D7F",
x"A1127D4E",
x"A0AC7D11",
x"A0327CB7",
x"9FA27C40",
x"9EF87BA3",
x"9E387AE5",
x"9D697A11",
x"9C977934",
x"9BD57865",
x"9B3577B9",
x"9AC97746",
x"9AA6771B",
x"9AD77740",
x"9B6677B9",
x"9C53787C",
x"9D9A797C",
x"9F317AA3",
x"A10A7BDE",
x"A3127D19",
x"A5387E44",
x"A76A7F56",
x"A996804F",
x"ABB1812F",
x"ADA981FD",
x"AF7B82BB",
x"B11B836B",
x"B281840F",
x"B3A6849E",
x"B487850D",
x"B51C854F",
x"B566855C",
x"B567852E",
x"B52884C2",
x"B4B38425",
x"B41C8366",
x"B377829C",
x"B2DC81E4",
x"B2608157",
x"B219810A",
x"B218810C",
x"B2668161",
x"B3048204",
x"B3EA82E3",
x"B50E83E8",
x"B65B84F7",
x"B7BC85F6",
x"B91686C8",
x"BA5A8760",
x"BB7487B3",
x"BC5E87C6",
x"BD1B87A7",
x"BDB2876C",
x"BE398731",
x"BEC78718",
x"BF74873E",
x"C05387B6",
x"C16D888B",
x"C2B489B5",
x"C40F8B1D",
x"C5498C94",
x"C61C8DE3",
x"C6358ECB",
x"C53F8F07",
x"C2EF8E60",
x"BF118CAC",
x"B98F89DA",
x"B28085FA",
x"AA218133",
x"A0D77BCE",
x"9729761F",
x"8DAA708A",
x"84ED6B6D",
x"7D75671D",
x"779D63D2",
x"739D61AB",
x"717660A8",
x"70FF60A8",
x"71E86176",
x"73CB62CF",
x"7637646C",
x"78C26609",
x"7B1B6772",
x"7D066886",
x"7E6A693A",
x"7F4E6991",
x"7FCE69A6",
x"80146997",
x"80526987",
x"80B16997",
x"815269DF",
x"82416A6B",
x"837C6B3A",
x"84F36C42",
x"868B6D6F",
x"88286EAB",
x"89AD6FDB",
x"8AFE70E8",
x"8C1371C5",
x"8CE57268",
x"8D7A72D2",
x"8DE07308",
x"8E247317",
x"8E59730C",
x"8E8A72F6",
x"8EC272E1",
x"8F0372D1",
x"8F4972C8",
x"8F8A72C0",
x"8FBB72AF",
x"8FC97285",
x"8FA97236",
x"8F4F71B4",
x"8EB470F8",
x"8DD77002",
x"8CC36EDB",
x"8B846D90",
x"8A2F6C37",
x"88DA6AEC",
x"87A169C8",
x"869768E3",
x"85CE684F",
x"85526814",
x"85246831",
x"853F689E",
x"85976948",
x"861A6A19",
x"86B56AF3",
x"87566BC4",
x"87EF6C75",
x"88776CF9",
x"88ED6D4F",
x"89556D76",
x"89BC6D7A",
x"8A2E6D69",
x"8AB96D4F",
x"8B676D3F",
x"8C3F6D44",
x"8D3E6D65",
x"8E596DA7",
x"8F816E06",
x"90A16E7D",
x"919F6F02",
x"92666F88",
x"92E07002",
x"93007066",
x"92C270A9",
x"922970C1",
x"914270AB",
x"90217065",
x"8EDF6FF0",
x"8D956F54",
x"8C626E97",
x"8B5C6DC5",
x"8A936CEF",
x"8A156C23",
x"89E66B70",
x"8A016AE9",
x"8A5F6A97",
x"8AF16A87",
x"8BAA6ABE",
x"8C776B3B",
x"8D4D6BFC",
x"8E226CF3",
x"8EEC6E12",
x"8FA76F45",
x"90527078",
x"90EE7195",
x"9180728A",
x"9207734A",
x"928573CB",
x"92FD740C",
x"936D7412",
x"93CF73E8",
x"9421739C",
x"945A733D",
x"947472DA",
x"9467727C",
x"942E722B",
x"93C371E9",
x"932871AF",
x"925F7175",
x"916F7133",
x"906470DF",
x"8F4C7076",
x"8E356FF6",
x"8D2A6F5E",
x"8C2E6EB5",
x"8B426E03",
x"8A5C6D4A",
x"896A6C90",
x"88556BD4",
x"87016B11",
x"855C6A45",
x"83586969",
x"80F9687A",
x"7E50677C",
x"7B896677",
x"78D8657F",
x"767F64A8",
x"74BF640B",
x"73D863C2",
x"73F363DD",
x"7525646C",
x"776B656C",
x"7A9E66D3",
x"7E8B6890",
x"82E86A8A",
x"87636CA4",
x"8BB66EC4",
x"8FA270D5",
x"92FE72C8",
x"95B97497",
x"97D97643",
x"997977D0",
x"9AC07946",
x"9BDF7AAD",
x"9D027C0C",
x"9E537D67",
x"9FEC7EBC",
x"A1DC800A",
x"A4268151",
x"A6C2828E",
x"A99E83C3",
x"ACA884F1",
x"AFC9861F",
x"B2F18753",
x"B6148895",
x"B92389EA",
x"BC1E8B53",
x"BEFC8CCE",
x"C1BC8E52",
x"C45A8FD6",
x"C6D0914C",
x"C91292A3",
x"CB1593CB",
x"CCC794B5",
x"CE199559",
x"CEFE95B1",
x"CF6895B8",
x"CF549576",
x"CEC794F2",
x"CDCD9435",
x"CC7A9351",
x"CAE79252",
x"C9339147",
x"C77C9039",
x"C5D98F34",
x"C45A8E39",
x"C3078D4C",
x"C1DB8C69",
x"C0D08B8A",
x"BFD68AAC",
x"BEDB89CC",
x"BDD788E7",
x"BCC48801",
x"BBA3871E",
x"BA818645",
x"B96B857E",
x"B87584D3",
x"B7B08447",
x"B72583DE",
x"B6D68397",
x"B6BF836D",
x"B6CF8359",
x"B6F58357",
x"B7208363",
x"B742837D",
x"B75383A8",
x"B75A83EE",
x"B767845D",
x"B79284FE",
x"B7F485E0",
x"B8A88704",
x"B9BF8867",
x"BB4289FE",
x"BD258BB2",
x"BF508D62",
x"C19F8EEC",
x"C3E19028",
x"C5E790F9",
x"C77E9145",
x"C88590FE",
x"C8E7902D",
x"C8A38EDD",
x"C7CA8D35",
x"C67E8B5C",
x"C4EA8983",
x"C34387D4",
x"C1B5867A",
x"C064858D",
x"BF678518",
x"BEC38514",
x"BE6A856D",
x"BE448601",
x"BE2F86AB",
x"BE0C8745",
x"BDC087B2",
x"BD4287E2",
x"BC9287D4",
x"BBC98799",
x"BB05874A",
x"BA6E870A",
x"BA2886F7",
x"BA4A8729",
x"BADC87AE",
x"BBCA887D",
x"BCF3897B",
x"BE1E8A85",
x"BF0A8B69",
x"BF7A8BF6",
x"BF3D8C06",
x"BE398B81",
x"BC688A62",
x"B9EB88BB",
x"B6F486B1",
x"B3C68474",
x"B0AC8239",
x"ADE38030",
x"AB997E7F",
x"A9DC7D32",
x"A89A7C43",
x"A7A87B99",
x"A6BF7B0B",
x"A5917A65",
x"A3D27979",
x"A1427823",
x"9DC0764B",
x"994D73F4",
x"940B7133",
x"8E3E6E33",
x"883E6B28",
x"82766852",
x"7D4665E8",
x"790A6418",
x"75FD6306",
x"744262B7",
x"73D96327",
x"74A76439",
x"767565C8",
x"790467A4",
x"7C1069A0",
x"7F566B90",
x"82A46D57",
x"85D86EE1",
x"88DC7027",
x"8BB2712E",
x"8E607208",
x"90F972C4",
x"938A7379",
x"9621743B",
x"98C67515",
x"9B79760C",
x"9E327725",
x"A0E67857",
x"A38A799C",
x"A60F7AEA",
x"A8717C34",
x"AAA97D77",
x"ACB97EAC",
x"AE9E7FD0",
x"B06080E8",
x"B1FE81F2",
x"B37882F1",
x"B4CA83E4",
x"B5F084CD",
x"B6DE85A7",
x"B794866C",
x"B8058719",
x"B83387A9",
x"B81F8817",
x"B7CD8862",
x"B747888A",
x"B6988894",
x"B5CA8885",
x"B4EB8867",
x"B407883F",
x"B3258817",
x"B24D87F1",
x"B18287D3",
x"B0C787BB",
x"B01B87A5",
x"AF7E878D",
x"AEED8769",
x"AE668733",
x"ADE686E9",
x"AD6E8683",
x"ACFF8605",
x"AC9C8571",
x"AC4784D0",
x"AC0B842C",
x"ABEE8391",
x"ABFA830A",
x"AC3582A2",
x"ACA68264",
x"AD4F8253",
x"AE2E8272",
x"AF3C82C2",
x"B06D833B",
x"B1B583D6",
x"B304848B",
x"B44D854F",
x"B5858618",
x"B6A886DC",
x"B7B58795",
x"B8B08840",
x"B9A388DA",
x"BA988966",
x"BB9689E4",
x"BCA68A59",
x"BDC98AC8",
x"BEFC8B32",
x"C0398B9E",
x"C1778C08",
x"C2AC8C76",
x"C3D08CE6",
x"C4E18D5B",
x"C5DD8DD6",
x"C6C48E5D",
x"C79F8EF1",
x"C8718F94",
x"C93A9042",
x"C9F990F7",
x"CAA991A8",
x"CB3E9249",
x"CBAA92CC",
x"CBDF9321",
x"CBD1933F",
x"CB7B9323",
x"CADE92CC",
x"CA059248",
x"C8FE91A7",
x"C7E19100",
x"C6C19065",
x"C5B58FE7",
x"C4C68F8E",
x"C3F88F55",
x"C3468F2C",
x"C2A08EFD",
x"C1F28EAC",
x"C12C8E1E",
x"C03A8D3E",
x"BF168C06",
x"BDC48A7D",
x"BC4D88B8",
x"BAC986DC",
x"B94C850F",
x"B7EB837A",
x"B6B08235",
x"B59B8150",
x"B49580C3",
x"B37B8074",
x"B21C8035",
x"B0427FD4",
x"ADBC7F19",
x"AA647DDA",
x"A6297BFB",
x"A11A7977",
x"9B607667",
x"953F72F9",
x"8F126F6B",
x"893B6C04",
x"841D6910",
x"800766C5",
x"7D35654F",
x"7BC164C1",
x"7BA16511",
x"7CB46624",
x"7EB567CC",
x"815D69D5",
x"845C6C07",
x"876C6E31",
x"8A597031",
x"8D0471F2",
x"8F69736B",
x"919474A1",
x"939E75A7",
x"95A8768F",
x"97D07768",
x"9A247841",
x"9CA77920",
x"9F497A06",
x"A1EE7AE8",
x"A4707BBD",
x"A6A67C74",
x"A8707D04",
x"A9B97D61",
x"AA7D7D8E",
x"AACC7D8B",
x"AAC27D65",
x"AA8A7D28",
x"AA547CE4",
x"AA4C7CA9",
x"AA957C84",
x"AB457C7C",
x"AC607C96",
x"ADD97CCD",
x"AF987D1E",
x"B17B7D7E",
x"B3577DE3",
x"B50B7E44",
x"B6757E9C",
x"B7827EEA",
x"B8297F2B",
x"B86D7F68",
x"B85A7FA6",
x"B8077FEE",
x"B78C8043",
x"B70280AC",
x"B6828128",
x"B61F81B7",
x"B5E58253",
x"B5DE82F7",
x"B60B8399",
x"B6648432",
x"B6DE84BB",
x"B768852E",
x"B7EE8584",
x"B85685BC",
x"B88A85CF",
x"B87485BC",
x"B8048581",
x"B7358519",
x"B6028488",
x"B47D83D0",
x"B2B682F7",
x"B0CC8204",
x"AEE08107",
x"AD17800C",
x"AB917F26",
x"AA677E64",
x"A9AB7DCF",
x"A9617D6D",
x"A9847D41",
x"AA047D46",
x"AAC77D6F",
x"ABB67DB2",
x"ACB57DFB",
x"ADA87E3D",
x"AE817E6E",
x"AF327E85",
x"AFB67E82",
x"B0087E6A",
x"B02E7E43",
x"B0267E19",
x"AFF77DF4",
x"AF9B7DD9",
x"AF127DC9",
x"AE577DBD",
x"AD637DAF",
x"AC2F7D8F",
x"AAB67D4E",
x"A8FA7CE3",
x"A6FF7C40",
x"A4D27B65",
x"A2807A57",
x"A01F7920",
x"9DC377D2",
x"9B837685",
x"9970754E",
x"979B7441",
x"960B736F",
x"94C272DC",
x"93B9728C",
x"92E47270",
x"9232727F",
x"919172A0",
x"90EE72C1",
x"904172CD",
x"8F7E72B1",
x"8EAA7266",
x"8DC671E8",
x"8CE5713A",
x"8C117066",
x"8B596F79",
x"8AC96E82",
x"8A606D90",
x"8A186CB0",
x"89DD6BE6",
x"89956B34",
x"891F6A94",
x"885569FA",
x"87146956",
x"85426896",
x"82CF67A5",
x"7FB86676",
x"7C0964FF",
x"77DC633E",
x"73596139",
x"6EAD5F01",
x"6A0A5CAC",
x"65A35A57",
x"61A1581F",
x"5E2A5621",
x"5B575477",
x"59335332",
x"57C3525D",
x"56FF51F7",
x"56D851F8",
x"573A5251",
x"580D52ED",
x"593753B3",
x"5AA1548F",
x"5C31556E",
x"5DD5563F",
x"5F7956FA",
x"610F5799",
x"6289581E",
x"63E2588C",
x"651258EB",
x"66145942",
x"66EE599A",
x"679E59F8",
x"682A5A64",
x"68995AE1",
x"68F35B6D",
x"69415C07",
x"69875CA8",
x"69CF5D49",
x"6A1D5DE3",
x"6A725E6C",
x"6ACE5EDD",
x"6B305F2F",
x"6B925F62",
x"6BEF5F73",
x"6C415F67",
x"6C805F46",
x"6CA75F15",
x"6CB15EE0",
x"6C9B5EAB",
x"6C685E7C",
x"6C175E57",
x"6BB25E3C",
x"6B3F5E2C",
x"6AC95E24",
x"6A5E5E24",
x"6A095E2C",
x"69D55E3D",
x"69CB5E5A",
x"69F25E87",
x"6A475EC3",
x"6AC95F11",
x"6B725F6D",
x"6C315FD3",
x"6CFD6039",
x"6DC7609A",
x"6E7F60E9",
x"6F1D6121",
x"6F9A613F",
x"6FF56142",
x"70306131",
x"70526110",
x"706860E9",
x"707960C6",
x"708F60B1",
x"70B160A9",
x"70DF60B2",
x"711960C9",
x"715560E6",
x"71896103",
x"71AA6115",
x"71AD6118",
x"71876108",
x"713860E7",
x"70BE60BB",
x"70246088",
x"6F75605C",
x"6EC5603E",
x"6E256038",
x"6DAA604D",
x"6D636080",
x"6D5C60CB",
x"6D9A6124",
x"6E1B6183",
x"6ED961DA",
x"6FC2621F",
x"70C86249",
x"71D66253",
x"72D8623E",
x"73BB620E",
x"747261CC",
x"74F06183",
x"7532613C",
x"75356100",
x"750060D2",
x"749760B4",
x"7409609E",
x"7362608B",
x"72B26070",
x"72076043",
x"716F5FFD",
x"70F35F9E",
x"70975F27",
x"705E5E9F",
x"70425E15",
x"703B5D95",
x"703A5D2B",
x"70315CE1",
x"70145CBF",
x"6FD45CC1",
x"6F6B5CE3",
x"6ED55D1B",
x"6E195D5C",
x"6D3E5D9A",
x"6C525DCC",
x"6B665DEA",
x"6A865DF3",
x"69C15DE7",
x"691B5DC9",
x"68965D9F",
x"682A5D6C",
x"67CC5D31",
x"676C5CEC",
x"66F85C95",
x"665B5C29",
x"65895B9F",
x"64785AF1",
x"63265A1C",
x"61995922",
x"5FDB580C",
x"5DFD56E6",
x"5C1955BF",
x"5A4154AB",
x"589053BA",
x"571952FE",
x"55EB527E",
x"5512523F",
x"5493523D",
x"546B5272",
x"549552D1",
x"55055349",
x"55B153C9",
x"568A5443",
x"578354AF",
x"588F5502",
x"59A6553F",
x"5ABE5568",
x"5BD55588",
x"5CE955A8",
x"5DF855D3",
x"5F005615",
x"60035674",
x"60FD56F4",
x"61EE5795",
x"62CE584F",
x"6399591A",
x"644A59EA",
x"64DB5AB3",
x"65495B6A",
x"65995C07",
x"65C95C82",
x"65E35CDF",
x"65F35D1C",
x"66045D43",
x"66215D5C",
x"66545D6D",
x"66A05D7E",
x"67075D95",
x"67825DB2",
x"68075DD3",
x"68875DF1",
x"68F25E08",
x"693A5E10",
x"69555E01",
x"69405DDA",
x"68FC5D9A",
x"68995D43",
x"68265CDF",
x"67B85C76",
x"676B5C14",
x"674F5BC8",
x"67755B9B",
x"67E35B98",
x"68995BC2",
x"69895C1A",
x"6AA15C9C",
x"6BCC5D41",
x"6CEF5DF8",
x"6DF35EB8",
x"6EC85F6E",
x"6F63600E",
x"6FC2608B",
x"6FEC60DF",
x"6FED6107",
x"6FD86107",
x"6FBE60E4",
x"6FAE60AD",
x"6FB4606D",
x"6FD86033",
x"7016600D",
x"70686004",
x"70C1601F",
x"7117605F",
x"715B60C1",
x"7183613C",
x"718D61C8",
x"71766258",
x"714562DD",
x"7103634F",
x"70BB63A1",
x"707563CF",
x"703863D3",
x"700963AF",
x"6FE36368",
x"6FC56301",
x"6FA56287",
x"6F7C6203",
x"6F446180",
x"6EFA6107",
x"6E9E60A1",
x"6E386052",
x"6DCF601D",
x"6D6E6001",
x"6D1E5FFC",
x"6CEB6006",
x"6CD6601A",
x"6CE36032",
x"6D0D6048",
x"6D4F6056",
x"6DA1605C",
x"6DF96059",
x"6E51604C",
x"6EA06039",
x"6EE56022",
x"6F1A600A",
x"6F425FF0",
x"6F595FD8",
x"6F5F5FBF",
x"6F545FA8",
x"6F315F92",
x"6EF95F7C",
x"6EAA5F64",
x"6E415F4C",
x"6DC25F35",
x"6D315F1E",
x"6C915F07",
x"6BE85EED",
x"6B3A5ECF",
x"6A895EA8",
x"69D55E73",
x"69195E29",
x"684F5DC6",
x"67755D46",
x"66865CA7",
x"657F5BEA",
x"64665B17",
x"63455A35",
x"62285952",
x"6123587D",
x"604757C5",
x"5FA6573C",
x"5F4E56ED",
x"5F4556E6",
x"5F8D5726",
x"602157B3",
x"60F65884",
x"61FF598E",
x"63315AC3",
x"64805C10",
x"65E85D62",
x"67665EA7",
x"68FD5FD0",
x"6AB060D5",
x"6C8261AD",
x"6E756259",
x"708662E0",
x"72B16350",
x"74EF63B8",
x"77346428",
x"797764B2",
x"7BB56566",
x"7DE8664C",
x"8011676C",
x"823468C1",
x"84586A42",
x"867D6BE1",
x"88A56D89",
x"8ACB6F23",
x"8CE37099",
x"8EDD71D8",
x"90A772D1",
x"922B737B",
x"935973D4",
x"942673E4",
x"948D73B7",
x"9492735F",
x"944372F2",
x"93B47282",
x"92FA7223",
x"922E71E5",
x"916671D2",
x"90B471EE",
x"90257236",
x"8FC372A1",
x"8F917326",
x"8F9173B4",
x"8FC1743D",
x"901E74B3",
x"90A47508",
x"914F7536",
x"9218753B",
x"92F47517",
x"93D774D2",
x"94B67474",
x"95817405",
x"96287393",
x"96A27327",
x"96E772C8",
x"96F4727C",
x"96D07244",
x"96847220",
x"961C720D",
x"95A97209",
x"953B7210",
x"94DD7223",
x"94977240",
x"946F7268",
x"9463729D",
x"947372E4",
x"949A733E",
x"94D273AC",
x"951A742A",
x"956D74B9",
x"95C9754D",
x"962B75DE",
x"968B7665",
x"96E376D7",
x"9725772C",
x"9743775E",
x"9731776F",
x"96DF775E",
x"96497734",
x"956E76F7",
x"945676AF",
x"93127664",
x"91BC761A",
x"906D75D4",
x"8F41758F",
x"8E507546",
x"8DAB74F1",
x"8D57748B",
x"8D52740F",
x"8D8B737C",
x"8DF172D8",
x"8E6D722F",
x"8EE9718C",
x"8F557103",
x"8FA970A6",
x"8FE77082",
x"901A70A1",
x"904F7108",
x"909A71B0",
x"910B7290",
x"91B4739A",
x"929474BA",
x"93AC75DB",
x"94ED76EE",
x"964377E4",
x"979778AF",
x"98CA794D",
x"99C979B9",
x"9A8379F5",
x"9AED7A05",
x"9B0879ED",
x"9AE079B3",
x"9A80795B",
x"99FB78EB",
x"995F7865",
x"98B477CA",
x"97F9771C",
x"971F7654",
x"96127571",
x"94B47468",
x"92E07334",
x"907D71CB",
x"8D74702B",
x"89C56E55",
x"857F6C4E",
x"80C86A27",
x"7BDB67F6",
x"770165DC",
x"728C63F9",
x"6EC7626C",
x"6BF86155",
x"6A4B60C5",
x"69D960C6",
x"6A9A6150",
x"6C6B6252",
x"6F1663AD",
x"7251653B",
x"75CE66D6",
x"7947685E",
x"7C7C69B1",
x"7F426AC1",
x"81866B89",
x"83466C0F",
x"84976C61",
x"85986C96",
x"86716CC1",
x"87466CF9",
x"88386D4A",
x"895C6DBD",
x"8AB96E4F",
x"8C4F6F00",
x"8E126FC4",
x"8FEE7094",
x"91D27168",
x"93A8723A",
x"95627309",
x"96F373D2",
x"98547496",
x"99847555",
x"9A80760D",
x"9B4876B9",
x"9BDC7750",
x"9C3C77CB",
x"9C697826",
x"9C61785B",
x"9C29786E",
x"9BC97865",
x"9B46784B",
x"9AAE782F",
x"9A0B781D",
x"996A7820",
x"98D4783E",
x"984F7877",
x"97D878C0",
x"976C790B",
x"97047948",
x"96957968",
x"9617795D",
x"9581791F",
x"94D578B2",
x"9414781D",
x"93467771",
x"927B76BD",
x"91C07616",
x"9127758B",
x"90B87523",
x"908074E5",
x"908074CB",
x"90B474D1",
x"911474E8",
x"9194750B",
x"9224752D",
x"92B4754E",
x"9335756A",
x"939B7585",
x"93DF75A3",
x"93FA75CA",
x"93F375FC",
x"93CD763D",
x"9397768C",
x"936276E7",
x"9342774A",
x"934977B3",
x"938D7820",
x"941A7890",
x"94F77902",
x"96257977",
x"979879ED",
x"99397A5E",
x"9AEA7AC9",
x"9C877B1F",
x"9DE77B5A",
x"9EEA7B6B",
x"9F6E7B4A",
x"9F667AF1",
x"9ECC7A60",
x"9DAB799B",
x"9C1C78B0",
x"9A4A77B0",
x"985F76B1",
x"968B75CA",
x"94FE750F",
x"93DA748D",
x"93387450",
x"93227458",
x"939074A0",
x"946D751C",
x"959A75BA",
x"96EE766A",
x"98437715",
x"997177AA",
x"9A5A781C",
x"9AE97860",
x"9B0E7872",
x"9ACC7850",
x"9A297801",
x"9936778B",
x"980776F9",
x"96B2765B",
x"954F75BE",
x"93F3752F",
x"92B174B9",
x"91957465",
x"90A9743A",
x"8FF37436",
x"8F6C744E",
x"8F077476",
x"8EB1749A",
x"8E4974A0",
x"8DAE746C",
x"8CB873E4",
x"8B3E72F1",
x"89217182",
x"864C6F93",
x"82BC6D2A",
x"7E866A5C",
x"79D1674B",
x"74DE6424",
x"6FF96118",
x"6B7A5E5D",
x"67BA5C25",
x"64FF5A94",
x"638359C5",
x"636259C0",
x"64995A7B",
x"67075BDD",
x"6A765DC2",
x"6E975FF7",
x"73186250",
x"77AB649E",
x"7C0766BC",
x"7FFC6894",
x"836D6A1D",
x"86566B59",
x"88C96C5B",
x"8AE26D38",
x"8CC56E0A",
x"8E956EEB",
x"90736FEB",
x"92707117",
x"94907272",
x"96CD73F2",
x"99147588",
x"9B4D771F",
x"9D5C789F",
x"9F2B79F4",
x"A0A57B06",
x"A1C67BCE",
x"A2907C46",
x"A30E7C71",
x"A3577C5E",
x"A3857C23",
x"A3B37BD9",
x"A3FB7B9B",
x"A4697B81",
x"A5047BA0",
x"A5C27BFE",
x"A68D7C99",
x"A7437D60",
x"A7BD7E35",
x"A7CF7EF1",
x"A7547F6D",
x"A6357F87",
x"A4677F1F",
x"A1F87E2D",
x"9F087CB4",
x"9BC87ACD",
x"9874789F",
x"954D7660",
x"928D7440",
x"905D7274",
x"8ED5711F",
x"8DF47051",
x"8DA5700D",
x"8DC1703D",
x"8E1170C0",
x"8E63716E",
x"8E877219",
x"8E5A72A1",
x"8DCF72EF",
x"8CE572FC",
x"8BB172CD",
x"8A527275",
x"88ED7212",
x"87A571BA",
x"86987186",
x"85D67180",
x"856571A9",
x"853A71F2",
x"853F7245",
x"855B7288",
x"856D729A",
x"855F726B",
x"851A71E9",
x"84947119",
x"83D37008",
x"82E96ECD",
x"81F06D8F",
x"81106C73",
x"80746BA1",
x"804B6B3D",
x"80BB6B5B",
x"81E36C0A",
x"83D26D48",
x"86886F05",
x"89F47126",
x"8DF17388",
x"924C75FF",
x"96C87862",
x"9B217A8C",
x"9F187C59",
x"A2777DB2",
x"A5127E8B",
x"A6D07EE3",
x"A7AB7EC6",
x"A7AF7E46",
x"A6F57D7F",
x"A5A87C8F",
x"A3F77B93",
x"A2177AA6",
x"A03979DD",
x"9E8A7946",
x"9D2878E2",
x"9C2978B4",
x"9B9278AF",
x"9B5A78C4",
x"9B6B78E2",
x"9BA978F9",
x"9BED78F9",
x"9C1778D6",
x"9C07788B",
x"9BA87816",
x"9AF1777B",
x"99E376C1",
x"988E75F2",
x"97037517",
x"955A7439",
x"93A7735B",
x"91F1727E",
x"903971A0",
x"8E7170B9",
x"8C806FBE",
x"8A486EA9",
x"87AC6D6E",
x"84976C07",
x"81006A73",
x"7CF368B7",
x"788D66DB",
x"740364EC",
x"6F9162FD",
x"6B7F6122",
x"680C5F70",
x"65705DF8",
x"63D25CCC",
x"63425BF6",
x"63BA5B7B",
x"651C5B5F",
x"673E5B9F",
x"69EC5C33",
x"6CEF5D12",
x"70175E32",
x"733A5F81",
x"763E60F4",
x"7916627E",
x"7BBF6411",
x"7E4565A4",
x"80B4672E",
x"831D68AD",
x"85906A1C",
x"88156B7C",
x"8AB56CCF",
x"8D6A6E19",
x"902E6F5B",
x"92F07097",
x"95A171CF",
x"98297303",
x"9A7A742C",
x"9C7E7547",
x"9E2E7650",
x"9F80773D",
x"A079780C",
x"A12478BA",
x"A1927948",
x"A1DD79B7",
x"A21E7A0C",
x"A2707A4E",
x"A2E97A84",
x"A3977AB4",
x"A4807AE4",
x"A59B7B18",
x"A6D77B51",
x"A8197B8F",
x"A9437BCE",
x"AA367C0C",
x"AAD97C43",
x"AB177C6F",
x"AAED7C8C",
x"AA637C96",
x"A9887C8F",
x"A87D7C78",
x"A75D7C53",
x"A64A7C25",
x"A5607BF2",
x"A4B27BC0",
x"A44C7B91",
x"A4297B65",
x"A4437B3D",
x"A4887B12",
x"A4E47AE1",
x"A5427AA2",
x"A5917A51",
x"A5C379EB",
x"A5D27972",
x"A5BF78EF",
x"A58D786A",
x"A54977F2",
x"A4FE7799",
x"A4BC776E",
x"A492777E",
x"A48E77CE",
x"A4B87861",
x"A518792D",
x"A5AE7A25",
x"A6787B34",
x"A76E7C46",
x"A8827D41",
x"A9A57E19",
x"AAC27EBD",
x"ABC57F2C",
x"AC9F7F68",
x"AD3F7F7B",
x"AD9F7F72",
x"ADBC7F5E",
x"AD987F4C",
x"AD3C7F43",
x"ACB87F4D",
x"AC187F68",
x"AB6E7F8F",
x"AAC97FB9",
x"AA307FDB",
x"A9AC7FEE",
x"A9387FEA",
x"A8CF7FCD",
x"A8667F99",
x"A7F37F50",
x"A7667EFC",
x"A6B87EA0",
x"A5DE7E46",
x"A4D77DED",
x"A3A87D98",
x"A2577D43",
x"A0F37CEA",
x"9F8B7C85",
x"9E337C11",
x"9CFD7B86",
x"9BF67AE7",
x"9B2B7A33",
x"9A9F7971",
x"9A5278A5",
x"9A3B77D8",
x"9A4C7712",
x"9A747657",
x"9A9C75AC",
x"9AB1750F",
x"9A987480",
x"9A4273FC",
x"999A7378",
x"989472EE",
x"97257254",
x"954B71A1",
x"930570CF",
x"905A6FD7",
x"8D5C6EB5",
x"8A1E6D6F",
x"86C36C0A",
x"836F6A94",
x"804F6924",
x"7D9467D1",
x"7B6D66B8",
x"7A0465F6",
x"797D65A5",
x"79E965D9",
x"7B4C6697",
x"7D9B67DE",
x"80B7699D",
x"84746BBA",
x"889E6E12",
x"8CFD7080",
x"915C72E5",
x"958E7525",
x"9976772F",
x"9D067902",
x"A0457AAA",
x"A3467C3F",
x"A62F7DDB",
x"A9297F99",
x"AC608198",
x"AFF883E3",
x"B40B867A",
x"B8A18955",
x"BDA98C58",
x"C3048F60",
x"C87E9244",
x"CDD494D8",
x"D2C696F9",
x"D70C988C",
x"DA749980",
x"DCD799D8",
x"DE26999D",
x"DE6E98EC",
x"DDD297E9",
x"DC8B96BD",
x"DADE9593",
x"D91A9497",
x"D78D93ED",
x"D67893AE",
x"D60C93EA",
x"D66494A1",
x"D78395C7",
x"D9559744",
x"DBB398F3",
x"DE619AAB",
x"E11D9C42",
x"E3A99D92",
x"E5C79E7B",
x"E7479EEC",
x"E80C9EE5",
x"E80D9E73",
x"E7579DB1",
x"E6009CC5",
x"E4379BD5",
x"E2299B07",
x"E0099A76",
x"DE039A33",
x"DC3D9A3B",
x"DACB9A80",
x"D9BA9AE6",
x"D9089B4A",
x"D8A79B87",
x"D8859B86",
x"D8899B33",
x"D89A9A89",
x"D8A69996",
x"D8989873",
x"D862973F",
x"D801961E",
x"D76C952E",
x"D6AA9487",
x"D5BE9434",
x"D4B39433",
x"D3959474",
x"D27494E5",
x"D15F9569",
x"D06A95E5",
x"CF9D963F",
x"CF069668",
x"CEA69655",
x"CE7B9603",
x"CE78957A",
x"CE8C94C4",
x"CEA393EC",
x"CEA59303",
x"CE7C9213",
x"CE189128",
x"CD6B9048",
x"CC748F76",
x"CB368EB1",
x"C9BC8DF7",
x"C8128D46",
x"C6508C97",
x"C4858BEA",
x"C2C68B39",
x"C1218A88",
x"BFA389D5",
x"BE598924",
x"BD468877",
x"BC7387D6",
x"BBE18740",
x"BB9386BD",
x"BB89864D",
x"BBC385F1",
x"BC4085AF",
x"BCFE8588",
x"BDFB8584",
x"BF3385A9",
x"C09F8604",
x"C239869E",
x"C3F7877D",
x"C5CE88A9",
x"C7B08A1F",
x"C9928BD9",
x"CB638DC8",
x"CD1B8FD5",
x"CEAD91EA",
x"D01693EA",
x"D15095BB",
x"D2549745",
x"D31C9873",
x"D3989934",
x"D3B0997C",
x"D3439940",
x"D2209872",
x"D0169709",
x"CCEE94F5",
x"C877922E",
x"C2918EAC",
x"BB358A76",
x"B27D8598",
x"A8A68036",
x"9E127A81",
x"933F74B4",
x"88BC6F1E",
x"7F1B6A09",
x"76E265BA",
x"7077626A",
x"6C19603E",
x"69D45F3B",
x"69895F53",
x"6AEB605C",
x"6D91621B",
x"7104644F",
x"74CF66B4",
x"78906910",
x"7C006B3A",
x"7EFC6D1A",
x"81836EAB",
x"83B16FF9",
x"85B27119",
x"87BB7221",
x"89FA732D",
x"8C8D744A",
x"8F7D757B",
x"92BE76BC",
x"962F77FE",
x"99A77930",
x"9CF37A3D",
x"9FE97B16",
x"A2667BB2",
x"A45A7C12",
x"A5C27C3D",
x"A6A87C46",
x"A7227C3D",
x"A74C7C3A",
x"A7407C4C",
x"A7157C7E",
x"A6DD7CD4",
x"A6A27D49",
x"A66A7DD1",
x"A6387E5D",
x"A60A7EDA",
x"A5E47F35",
x"A5C67F61",
x"A5B37F56",
x"A5AF7F0E",
x"A5B97E8F",
x"A5D27DE3",
x"A5F47D18",
x"A6187C40",
x"A6357B6F",
x"A6427AB7",
x"A6337A28",
x"A60579CA",
x"A5B579A5",
x"A54279B4",
x"A4B179F5",
x"A4057A5A",
x"A3467AD1",
x"A2767B4D",
x"A1987BB7",
x"A0AC7C02",
x"9FAF7C1F",
x"9EA17C04",
x"9D7B7BAC",
x"9C437B1C",
x"9AFD7A58",
x"99AF7971",
x"98677872",
x"9735776F",
x"9628767C",
x"955275A9",
x"94C17506",
x"947D749F",
x"948D747C",
x"94EC749D",
x"95927502",
x"967675A2",
x"9781766E",
x"98A47758",
x"99C6784B",
x"9AD77934",
x"9BC37A01",
x"9C7E7A9D",
x"9CFD7AFE",
x"9D3B7B19",
x"9D367AED",
x"9CF37A7B",
x"9C7879CE",
x"9BCF78F4",
x"9B0377FC",
x"9A1F76FB",
x"99327602",
x"98427521",
x"975C7467",
x"968373D7",
x"95BC7376",
x"95087340",
x"9467732F",
x"93D97339",
x"935A7357",
x"92ED7380",
x"929373B1",
x"924C73E4",
x"92217419",
x"9215744E",
x"922B7486",
x"926674BE",
x"92C074F2",
x"9335751C",
x"93B57534",
x"942F7534",
x"94927513",
x"94C974CD",
x"94C8745F",
x"948373CD",
x"93FA731D",
x"93367258",
x"92437188",
x"912F70B3",
x"900D6FDE",
x"8EE46F09",
x"8DB86E2D",
x"8C816D42",
x"8B316C3D",
x"89AE6B10",
x"87E269B7",
x"85B8682D",
x"83286679",
x"803864AD",
x"7CFD62DD",
x"79A06125",
x"76565FA2",
x"735B5E73",
x"70E65DAB",
x"6F2A5D59",
x"6E475D81",
x"6E445E1C",
x"6F165F18",
x"709B605C",
x"72A761CB",
x"74FF6345",
x"776D64AE",
x"79C765F0",
x"7BEA66FC",
x"7DCB67CF",
x"7F69686C",
x"80D668E1",
x"822A693F",
x"8379699C",
x"84DD6A09",
x"86626A9C",
x"880D6B5C",
x"89DA6C51",
x"8BBE6D75",
x"8DAB6EBD",
x"8F94701A",
x"916C7179",
x"932B72C7",
x"94D273F4",
x"965D74F2",
x"97CF75BC",
x"99277651",
x"9A5F76B4",
x"9B6E76F1",
x"9C4B770D",
x"9CE97716",
x"9D3F7712",
x"9D467708",
x"9D0176F9",
x"9C7B76E7",
x"9BC376CD",
x"9AF176A9",
x"9A1C767B",
x"995D7640",
x"98C375FB",
x"985D75B1",
x"982C756B",
x"982E752D",
x"985A7501",
x"98A774EC",
x"990A74F6",
x"997B751D",
x"99FB7562",
x"9A8A75C3",
x"9B2E7639",
x"9BEE76BD",
x"9CCF774B",
x"9DD077E0",
x"9EEE7877",
x"A01C790E",
x"A14C79A5",
x"A2667A3C",
x"A3577AD1",
x"A40E7B61",
x"A47A7BE8",
x"A4927C5B",
x"A4567CB3",
x"A3CA7CE3",
x"A2F87CDE",
x"A1EE7C9E",
x"A0B87C1E",
x"9F637B5E",
x"9DFE7A68",
x"9C927948",
x"9B297812",
x"99CF76DA",
x"988D75B3",
x"976C74B3",
x"967773E5",
x"95BC7354",
x"95437300",
x"951272E6",
x"952972FF",
x"9586733E",
x"961B7397",
x"96DA7403",
x"97AE7475",
x"987E74E7",
x"99387555",
x"99C675BA",
x"9A1A7613",
x"9A29765B",
x"99F3768F",
x"997A76A9",
x"98C976A6",
x"97ED7682",
x"96F8763E",
x"960075DC",
x"95177562",
x"945274DB",
x"93C37450",
x"937973CE",
x"937A7361",
x"93CB7312",
x"946372E8",
x"953472E5",
x"96257305",
x"971D7341",
x"97F97392",
x"989B73EA",
x"98E7743A",
x"98CF7479",
x"984C749C",
x"9763749A",
x"962B7471",
x"94BE741C",
x"933E739F",
x"91C97300",
x"907C724A",
x"8F627182",
x"8E7C70B4",
x"8DBB6FE9",
x"8D036F27",
x"8C2F6E6F",
x"8B1A6DBF",
x"89A16D10",
x"87AC6C57",
x"85356B89",
x"82486A9A",
x"7F006989",
x"7B8C6854",
x"78266703",
x"750C65AB",
x"72776463",
x"709D634C",
x"6FA16280",
x"6F96621B",
x"7079622D",
x"723A62BC",
x"74B563C1",
x"77C16524",
x"7B2866C8",
x"7EBC6889",
x"824F6A44",
x"85BE6BDB",
x"88EF6D3B",
x"8BD86E61",
x"8E766F55",
x"90D0702B",
x"92F770FF",
x"94FE71EB",
x"96F77305",
x"98F4745A",
x"9B0475EA",
x"9D3277AD",
x"9F80798E",
x"A1ED7B71",
x"A4717D3F",
x"A7037EE0",
x"A9918046",
x"AC0C8170",
x"AE5E8261",
x"B0778325",
x"B24283C9",
x"B3AD845A",
x"B4AF84DE",
x"B53F8557",
x"B55B85BD",
x"B5098605",
x"B4548621",
x"B3498607",
x"B1FB85AE",
x"B07E8519",
x"AEE18450",
x"AD368364",
x"AB878268",
x"A9DA8170",
x"A838808A",
x"A6A47FC3",
x"A5257F1E",
x"A3C27E99",
x"A2887E2C",
x"A1877DD3",
x"A0D07D85",
x"A0717D44",
x"A0797D16",
x"A0EB7D01",
x"A1C37D12",
x"A2F07D53",
x"A4527DC7",
x"A5C27E6B",
x"A7157F2F",
x"A81F8000",
x"A8B980BF",
x"A8CA814A",
x"A84C818A",
x"A749816A",
x"A5E180EA",
x"A4478015",
x"A2B87F0A",
x"A1707DEF",
x"A0AB7CF5",
x"A0957C47",
x"A1487C0B",
x"A2C27C57",
x"A4ED7D2D",
x"A7997E7B",
x"AA87801E",
x"AD6E81E6",
x"B00B839F",
x"B21E8517",
x"B37B8625",
x"B40E86B2",
x"B3DA86B9",
x"B2F58645",
x"B18C8570",
x"AFD3845E",
x"AE018338",
x"AC4A821C",
x"AAD48126",
x"A9BD8067",
x"A90E7FE0",
x"A8C37F8B",
x"A8D17F5B",
x"A9257F42",
x"A9A67F35",
x"AA427F29",
x"AAE87F1E",
x"AB8C7F16",
x"AC287F1C",
x"ACB37F33",
x"AD2C7F64",
x"AD8F7FAF",
x"ADD9800F",
x"ADFF807B",
x"AE0180E1",
x"ADD78136",
x"AD818167",
x"AD01816D",
x"AC548142",
x"AB8580E7",
x"AA998066",
x"A9987FC9",
x"A8877F1F",
x"A76D7E78",
x"A64A7DD9",
x"A5237D47",
x"A3F87CC3",
x"A2C57C44",
x"A1887BC0",
x"A0387B25",
x"9EC97A63",
x"9D297968",
x"9B407826",
x"98F77692",
x"962F74A5",
x"92D3725E",
x"8ED66FC1",
x"8A3B6CDE",
x"851469C4",
x"7F8E6690",
x"79E86362",
x"746C605F",
x"6F705DAE",
x"6B445B73",
x"682B59CA",
x"665658CA",
x"65D7587D",
x"66A058DC",
x"688A59D9",
x"6B595B56",
x"6EC55D32",
x"727F5F43",
x"76446164",
x"79E06376",
x"7D32655F",
x"802B6713",
x"82D2688E",
x"853269D8",
x"87656AFC",
x"897D6C0A",
x"8B8A6D12",
x"8D946E1E",
x"8F9A6F37",
x"919A705E",
x"938E7193",
x"957472D2",
x"974D7417",
x"9922755E",
x"9B0076A5",
x"9CF477EF",
x"9F0B793E",
x"A14F7A96",
x"A3BB7BF8",
x"A6437D63",
x"A8D47ED1",
x"AB4F803A",
x"AD94818F",
x"AF8882C3",
x"B11283C6",
x"B225848B",
x"B2BD850B",
x"B2E88545",
x"B2B6853C",
x"B24084FD",
x"B1A38497",
x"B0F48418",
x"B0478394",
x"AFA88315",
x"AF1582A6",
x"AE8A824A",
x"ADFE8201",
x"AD6681C6",
x"ACB88194",
x"ABEE8164",
x"AB0C8135",
x"AA198104",
x"A92480D1",
x"A83C80A6",
x"A7738082",
x"A6D3806D",
x"A6668064",
x"A628806A",
x"A6118075",
x"A60D807C",
x"A6078078",
x"A5ED805A",
x"A5AE801C",
x"A5427FBA",
x"A4AF7F37",
x"A4047E9E",
x"A35D7DFA",
x"A2DD7D5E",
x"A2A57CE0",
x"A2D37C91",
x"A37A7C7C",
x"A49B7CA9",
x"A6267D15",
x"A7FB7DB5",
x"A9EB7E74",
x"ABC27F3C",
x"AD4A7FF5",
x"AE5D808A",
x"AEDE80E8",
x"AEC98108",
x"AE2B80E8",
x"AD258091",
x"ABE6800F",
x"AA9C7F78",
x"A97A7EE0",
x"A8A27E51",
x"A8267DDA",
x"A8087D7C",
x"A8367D37",
x"A8917CFF",
x"A8F47CCD",
x"A9387C95",
x"A93F7C50",
x"A8F87BFE",
x"A8647BA6",
x"A7957B54",
x"A6AB7B1B",
x"A5CC7B09",
x"A5297B32",
x"A4EC7B9F",
x"A5367C54",
x"A61C7D4C",
x"A7A17E7A",
x"A9B97FC7",
x"AC4A8123",
x"AF2E8276",
x"B23B83AD",
x"B54684C0",
x"B82685AB",
x"BABD8671",
x"BCF4871B",
x"BEBF87B5",
x"C01B8845",
x"C10888D0",
x"C18B8955",
x"C1A289C5",
x"C1498A0D",
x"C0748A11",
x"BF0B89B5",
x"BCF488DA",
x"BA0E876D",
x"B63C855C",
x"B16B82A8",
x"AB957F5B",
x"A4C57B92",
x"9D1F776E",
x"94DD731D",
x"8C4F6ED1",
x"83CF6AB8",
x"7BC56701",
x"749663CF",
x"6E996139",
x"6A165F50",
x"673D5E15",
x"661A5D83",
x"66A65D8B",
x"68B45E1C",
x"6C095F21",
x"70556086",
x"75456237",
x"7A876421",
x"7FD26637",
x"84E96866",
x"89A16AA4",
x"8DE76CE3",
x"91B26F1D",
x"950D7143",
x"98077350",
x"9AB8753D",
x"9D357706",
x"9F8E78A9",
x"A1C97A22",
x"A3E67B71",
x"A5DC7C95",
x"A79B7D8C",
x"A9157E54",
x"AA397EED",
x"AB047F54",
x"AB727F91",
x"AB957FA6",
x"AB7E7F9F",
x"AB4C7F88",
x"AB1C7F71",
x"AB0E7F68",
x"AB367F7F",
x"ABA17FC0",
x"AC4D802D",
x"AD2C80CA",
x"AE28818A",
x"AF1F825E",
x"AFF18335",
x"B08083FA",
x"B0B38499",
x"B0828505",
x"AFEE8532",
x"AF05851E",
x"ADE084CD",
x"AC9B8449",
x"AB53839F",
x"AA2582E0",
x"A928821E",
x"A8698164",
x"A7EE80C3",
x"A7B98040",
x"A7BF7FE3",
x"A7F77FAD",
x"A8527F9E",
x"A8C57FB0",
x"A93F7FE1",
x"A9B88028",
x"AA22807A",
x"AA7480CF",
x"AAA58119",
x"AAAF8150",
x"AA8C8167",
x"AA3B8154",
x"A9BD8114",
x"A91A80A1",
x"A85A7FFB",
x"A78E7F2B",
x"A6C67E39",
x"A6117D2F",
x"A5807C1C",
x"A5197B0F",
x"A4E37A12",
x"A4D4792F",
x"A4E6786D",
x"A50177CB",
x"A512774D",
x"A50076EC",
x"A4B676A6",
x"A4297675",
x"A3527657",
x"A235764A",
x"A0E1764E",
x"9F6E7667",
x"9DF77695",
x"9C9576D8",
x"9B647733",
x"9A73779D",
x"99C67810",
x"995C7881",
x"992478E0",
x"99087922",
x"98F3793A",
x"98CD7925",
x"988A78E1",
x"98247877",
x"97A277F4",
x"971A776C",
x"969F76F7",
x"965276A5",
x"96487686",
x"969176A5",
x"973176FF",
x"98187789",
x"99347833",
x"9A5F78E4",
x"9B747985",
x"9C557A02",
x"9CE77A4A",
x"9D217A5B",
x"9D087A39",
x"9CB379EF",
x"9C407992",
x"9BD27934",
x"9B8378E7",
x"9B6478B0",
x"9B74788F",
x"9B9A7875",
x"9BAB784B",
x"9B7177F4",
x"9AAF7751",
x"992E764B",
x"96C874D2",
x"937072E6",
x"8F377097",
x"8A4C6E05",
x"84FB6B58",
x"7FA468C4",
x"7AA76679",
x"766964A4",
x"733B6365",
x"715262C9",
x"70CB62D5",
x"719E6376",
x"73A56493",
x"76A76609",
x"7A5867B4",
x"7E666972",
x"82866B27",
x"86716CC1",
x"89F76E37",
x"8CF16F85",
x"8F5370B0",
x"911E71BE",
x"926072BA",
x"933473A6",
x"93B97488",
x"94177561",
x"9470762D",
x"94E176EB",
x"95887796",
x"9671782D",
x"97A578B0",
x"991D791D",
x"9AC97979",
x"9C9279C6",
x"9E5A7A06",
x"9FFE7A3C",
x"A1607A68",
x"A2637A88",
x"A2F77A98",
x"A3127A95",
x"A2BB7A7B",
x"A2007A47",
x"A0FA79F8",
x"9FC8798E",
x"9E88790F",
x"9D5C787F",
x"9C5A77E5",
x"9B95774B",
x"9B1576B6",
x"9ADA762D",
x"9ADC75B7",
x"9B0D7557",
x"9B5C750C",
x"9BBB74D7",
x"9C1774B7",
x"9C6474A7",
x"9C9874A5",
x"9CAE74AD",
x"9C9F74B9",
x"9C6E74C6",
x"9C1A74CE",
x"9BA274D0",
x"9B0A74C6",
x"9A5074AF",
x"99777488",
x"98817451",
x"9770740D",
x"964873BB",
x"950B7362",
x"93C27300",
x"9271729C",
x"91247234",
x"8FE071CA",
x"8EAF715E",
x"8D9A70EB",
x"8CA47073",
x"8BD66FF3",
x"8B356F6F",
x"8AC16EE6",
x"8A7C6E62",
x"8A646DE5",
x"8A746D79",
x"8AA56D24",
x"8AEF6CE9",
x"8B456CCB",
x"8B9E6CC8",
x"8BEF6CD9",
x"8C2F6CFA",
x"8C596D21",
x"8C6A6D4A",
x"8C636D6E",
x"8C486D8A",
x"8C1D6DA0",
x"8BE96DB4",
x"8BB26DCB",
x"8B7D6DEB",
x"8B4C6E16",
x"8B216E51",
x"8AF96E9C",
x"8AD36EF3",
x"8AAE6F52",
x"8A896FB4",
x"8A647014",
x"8A43706E",
x"8A2E70BD",
x"8A277102",
x"8A32713D",
x"8A56716B",
x"8A90718F",
x"8ADC71A3",
x"8B3171A3",
x"8B81718C",
x"8BBE7155",
x"8BD970F9",
x"8BC67076",
x"8B7D6FCB",
x"8AFD6F00",
x"8A4B6E1C",
x"89746D28",
x"888A6C37",
x"879E6B4F",
x"86BC6A7C",
x"85ED69C1",
x"852E691B",
x"846D6881",
x"839167E5",
x"82796732",
x"80FD6658",
x"7EFA6544",
x"7C5E63EF",
x"79216255",
x"7556607E",
x"71275E80",
x"6CD25C71",
x"68A75A77",
x"64F858B5",
x"62175750",
x"60475666",
x"5FB3560B",
x"6068564D",
x"6258572B",
x"65585895",
x"692A5A77",
x"6D835CB1",
x"72165F22",
x"769E61A9",
x"7AE66427",
x"7EC96683",
x"823868AD",
x"85366A9C",
x"87D06C4D",
x"8A216DC8",
x"8C3E6F16",
x"8E437045",
x"90437161",
x"924F7275",
x"946D738D",
x"96A274AD",
x"98F375D7",
x"9B5A7709",
x"9DD3783E",
x"A053796D",
x"A2D07A89",
x"A5367B88",
x"A7707C5D",
x"A9677CFF",
x"AB027D67",
x"AC2D7D95",
x"ACDA7D8B",
x"AD017D53",
x"ACA87CFB",
x"ABDE7C94",
x"AABC7C30",
x"A9607BE3",
x"A7EA7BB4",
x"A67D7BB0",
x"A5337BD6",
x"A4257C1C",
x"A3607C78",
x"A2EB7CDB",
x"A2C77D35",
x"A2EE7D75",
x"A3537D96",
x"A3EC7D95",
x"A4A77D75",
x"A5767D41",
x"A6497D08",
x"A7127CD6",
x"A7C37CB9",
x"A8547CB6",
x"A8BC7CD0",
x"A8F57D02",
x"A9047D41",
x"A8E97D81",
x"A8AB7DB0",
x"A8537DC7",
x"A7E97DBC",
x"A7757D8F",
x"A6FE7D46",
x"A6877CED",
x"A6127C91",
x"A5A17C44",
x"A5367C13",
x"A4D47C09",
x"A4807C2D",
x"A43D7C7C",
x"A41A7CF4",
x"A4187D88",
x"A4427E2D",
x"A49C7ED7",
x"A5257F77",
x"A5D98005",
x"A6B0807A",
x"A79B80D3",
x"A88E8111",
x"A9778133",
x"AA4C8140",
x"AAFD813C",
x"AB858129",
x"ABDE810A",
x"AC0580DA",
x"ABF6809B",
x"ABAF8046",
x"AB2F7FD4",
x"AA747F40",
x"A97B7E85",
x"A8457D9F",
x"A6D67C8F",
x"A5367B5B",
x"A3707A0C",
x"A19778B0",
x"9FC07758",
x"9E037619",
x"9C787506",
x"9B387430",
x"9A5573A5",
x"99D9736E",
x"99CA738F",
x"9A267403",
x"9ADF74C3",
x"9BE175BA",
x"9D1176D7",
x"9E537801",
x"9F887922",
x"A0987A25",
x"A16A7AF5",
x"A1F47B8B",
x"A2337BDD",
x"A22B7BED",
x"A1EA7BC1",
x"A1817B65",
x"A1017AE3",
x"A07A7A46",
x"9FEE7995",
x"9F5978D4",
x"9EA777FE",
x"9DBC770D",
x"9C7475F4",
x"9AAA74A3",
x"983F7313",
x"951E713B",
x"91496F21",
x"8CD26CCE",
x"87E56A56",
x"82C167DB",
x"7DB16579",
x"79096358",
x"75176195",
x"7220604C",
x"70525F8E",
x"6FC65F60",
x"707A5FBE",
x"7253609D",
x"752061E6",
x"78A26383",
x"7C97655C",
x"80B96758",
x"84CF6962",
x"88A86B6C",
x"8C2A6D68",
x"8F4B6F4B",
x"92137114",
x"949872C0",
x"96F8744E",
x"995975C1",
x"9BD9771D",
x"9E92786B",
x"A19279AF",
x"A4D77AF1",
x"A8507C36",
x"ABDE7D81",
x"AF577ED4",
x"B28F8029",
x"B55A817E",
x"B79182CA",
x"B91F8404",
x"B9FC8521",
x"BA368619",
x"B9E786E7",
x"B9398785",
x"B85787F1",
x"B7728828",
x"B6AF882B",
x"B62587F9",
x"B5DB8794",
x"B5D086FE",
x"B5EA863C",
x"B60F8554",
x"B6228450",
x"B609833F",
x"B5B68232",
x"B529813C",
x"B46D8072",
x"B3997FE6",
x"B2CD7FA0",
x"B22B7FAB",
x"B1CA7FFE",
x"B1BF8091",
x"B20F814F",
x"B2B38222",
x"B39482F1",
x"B49283A5",
x"B58C8429",
x"B65D8471",
x"B6E58478",
x"B70F8442",
x"B6CD83D6",
x"B6238346",
x"B51B82A1",
x"B3CE81FB",
x"B25A8166",
x"B0E480ED",
x"AF8F809B",
x"AE828077",
x"ADD98080",
x"ADA980B5",
x"ADFF810E",
x"AEDE8187",
x"B03A8216",
x"B20082B5",
x"B411835A",
x"B64F8402",
x"B89484A8",
x"BAC2854A",
x"BCBD85E7",
x"BE748680",
x"BFDB8714",
x"C0F187A4",
x"C1B9882B",
x"C24088AB",
x"C291891E",
x"C2B6897E",
x"C2B989C9",
x"C29F89F7",
x"C2678A05",
x"C20E89EF",
x"C18B89B2",
x"C0D88952",
x"BFF188CD",
x"BED0882C",
x"BD7B8776",
x"BBF886AF",
x"BA5885E6",
x"B8AB8523",
x"B70A8473",
x"B58C83E1",
x"B44C8377",
x"B35E8340",
x"B2D4833F",
x"B2B38374",
x"B2FA83DD",
x"B39B8470",
x"B481851C",
x"B58C85D6",
x"B69F868A",
x"B7968729",
x"B85987AC",
x"B8D4880D",
x"B901884C",
x"B8E38870",
x"B8848880",
x"B7F58883",
x"B746887D",
x"B67F8867",
x"B59C8838",
x"B48F87DC",
x"B33D8736",
x"B17E862E",
x"AF2E84A9",
x"AC2B8299",
x"A8607FFC",
x"A3D07CE1",
x"9E947962",
x"98DD75AC",
x"92F471F4",
x"8D2E6E73",
x"87E06B5E",
x"836268DF",
x"7FF06717",
x"7DBA6611",
x"7CC965CB",
x"7D146630",
x"7E766721",
x"80B8687D",
x"839A6A20",
x"86DF6BE6",
x"8A4C6DB7",
x"8DB96F83",
x"910A7143",
x"943572F6",
x"973974A3",
x"9A267652",
x"9D0D780F",
x"A00079E0",
x"A30C7BC7",
x"A63F7DC7",
x"A9967FD9",
x"AD0E81F4",
x"B099840E",
x"B4298619",
x"B7A9880A",
x"BB0489D0",
x"BE258B66",
x"C0FB8CC3",
x"C3788DE5",
x"C5928ECC",
x"C7448F7C",
x"C88C8FFA",
x"C96E904E",
x"C9F1907A",
x"CA1F908A",
x"CA05907D",
x"C9B49056",
x"C93D9018",
x"C8B08FC2",
x"C81C8F51",
x"C7928EC8",
x"C71B8E2B",
x"C6BF8D80",
x"C6818CD0",
x"C6618C27",
x"C6578B91",
x"C65A8B1B",
x"C65E8AD0",
x"C6588AB5",
x"C6418ACD",
x"C6138B18",
x"C5D68B94",
x"C5948C3B",
x"C5608D06",
x"C5548DF4",
x"C5898F03",
x"C6199031",
x"C711917F",
x"C87792ED",
x"CA43947C",
x"CC619621",
x"CEB397D9",
x"D1199993",
x"D3719B40",
x"D5A09CD1",
x"D7989E3A",
x"D9549F71",
x"DADFA073",
x"DC4DA143",
x"DDB0A1E9",
x"DF1CA271",
x"E09CA2E4",
x"E22AA34A",
x"E3BAA3AA",
x"E530A3FF",
x"E668A447",
x"E745A474",
x"E7AEA47C",
x"E799A458",
x"E70AA404",
x"E61CA385",
x"E4F5A2E4",
x"E3C0A233",
x"E2ADA186",
x"E1E1A0EE",
x"E16CA078",
x"E14EA029",
x"E1719FFC",
x"E1A99FE1",
x"E1C19FBD",
x"E1809F73",
x"E0B09EE7",
x"DF2A9DF9",
x"DCE09C9C",
x"D9D39AC8",
x"D6259886",
x"D20695EC",
x"CDB7931A",
x"C97B903B",
x"C58F8D79",
x"C2298AFD",
x"BF6788E7",
x"BD53874F",
x"BBDB8636",
x"BADD8598",
x"BA268559",
x"B97A8557",
x"B8A1856A",
x"B7678567",
x"B5AF8527",
x"B36E848E",
x"B0B08391",
x"AD958230",
x"AA4D8080",
x"A70B7E9F",
x"A4057CB0",
x"A1647ADB",
x"9F3E7940",
x"9D8E77F1",
x"9C3F76F4",
x"9B1E763A",
x"99EF75A5",
x"986A750C",
x"96527443",
x"9373731F",
x"8FB37180",
x"8B176F5B",
x"85BE6CB3",
x"7FE569A6",
x"79DC665F");

begin
process(clka) 
begin 
	if(rising_edge(clka)) then
		if ena = '1' then
			douta <= ROM(to_integer(unsigned(addra (15 downto 0)))) ;
		end if;
	end if;
end process ;
end bijeibural;