----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:43:16 10/18/2016 
-- Design Name: 
-- Module Name:    mult_1bit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mult_1bit is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
			  pin : in  STD_LOGIC;
           cin : in  STD_LOGIC;
			  cout : out  STD_LOGIC;
           pout : out  STD_LOGIC);
           
end mult_1bit;

architecture Behavioral of mult_1bit is

begin
	pout <= (a and b) xor pin xor cin; 
	cout <= ((a and b) and pin) or (cin and ((a and b) xor pin));
end Behavioral;

